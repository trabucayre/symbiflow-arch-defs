`timescale 1ns/10ps
(* whitebox *)
module MULT (
	input [31:0] Amult,
	input [31:0] Bmult,
	input [1:0] Valid_mult,
	output [63:0] Cmult,
	input sel_mul_32x32
);

	(* DELAY_MATRIX_Amult="{iopath_Amult0_Cmult0} {iopath_Amult0_Cmult1} {iopath_Amult0_Cmult2} {iopath_Amult0_Cmult3} {iopath_Amult0_Cmult4} {iopath_Amult0_Cmult5} {iopath_Amult0_Cmult6} {iopath_Amult0_Cmult7} {iopath_Amult0_Cmult8} {iopath_Amult0_Cmult9} {iopath_Amult0_Cmult10} {iopath_Amult0_Cmult11} {iopath_Amult0_Cmult12} {iopath_Amult0_Cmult13} {iopath_Amult0_Cmult14} {iopath_Amult0_Cmult15} {iopath_Amult0_Cmult16} {iopath_Amult0_Cmult17} {iopath_Amult0_Cmult18} {iopath_Amult0_Cmult19} {iopath_Amult0_Cmult20} {iopath_Amult0_Cmult21} {iopath_Amult0_Cmult22} {iopath_Amult0_Cmult23} {iopath_Amult0_Cmult24} {iopath_Amult0_Cmult25} {iopath_Amult0_Cmult26} {iopath_Amult0_Cmult27} {iopath_Amult0_Cmult28} {iopath_Amult0_Cmult29} {iopath_Amult0_Cmult30} {iopath_Amult0_Cmult31} {iopath_Amult0_Cmult32} {iopath_Amult0_Cmult33} {iopath_Amult0_Cmult34} {iopath_Amult0_Cmult35} {iopath_Amult0_Cmult36} {iopath_Amult0_Cmult37} {iopath_Amult0_Cmult38} {iopath_Amult0_Cmult39} {iopath_Amult0_Cmult40} {iopath_Amult0_Cmult41} {iopath_Amult0_Cmult42} {iopath_Amult0_Cmult43} {iopath_Amult0_Cmult44} {iopath_Amult0_Cmult45} {iopath_Amult0_Cmult46} {iopath_Amult0_Cmult47} {iopath_Amult0_Cmult48} {iopath_Amult0_Cmult49} {iopath_Amult0_Cmult50} {iopath_Amult0_Cmult51} {iopath_Amult0_Cmult52} {iopath_Amult0_Cmult53} {iopath_Amult0_Cmult54} {iopath_Amult0_Cmult55} {iopath_Amult0_Cmult56} {iopath_Amult0_Cmult57} {iopath_Amult0_Cmult58} {iopath_Amult0_Cmult59} {iopath_Amult0_Cmult60} {iopath_Amult0_Cmult61} {iopath_Amult0_Cmult62} {iopath_Amult0_Cmult63} 0 {iopath_Amult1_Cmult1} {iopath_Amult1_Cmult2} {iopath_Amult1_Cmult3} {iopath_Amult1_Cmult4} {iopath_Amult1_Cmult5} {iopath_Amult1_Cmult6} {iopath_Amult1_Cmult7} {iopath_Amult1_Cmult8} {iopath_Amult1_Cmult9} {iopath_Amult1_Cmult10} {iopath_Amult1_Cmult11} {iopath_Amult1_Cmult12} {iopath_Amult1_Cmult13} {iopath_Amult1_Cmult14} {iopath_Amult1_Cmult15} {iopath_Amult1_Cmult16} {iopath_Amult1_Cmult17} {iopath_Amult1_Cmult18} {iopath_Amult1_Cmult19} {iopath_Amult1_Cmult20} {iopath_Amult1_Cmult21} {iopath_Amult1_Cmult22} {iopath_Amult1_Cmult23} {iopath_Amult1_Cmult24} {iopath_Amult1_Cmult25} {iopath_Amult1_Cmult26} {iopath_Amult1_Cmult27} {iopath_Amult1_Cmult28} {iopath_Amult1_Cmult29} {iopath_Amult1_Cmult30} {iopath_Amult1_Cmult31} {iopath_Amult1_Cmult32} {iopath_Amult1_Cmult33} {iopath_Amult1_Cmult34} {iopath_Amult1_Cmult35} {iopath_Amult1_Cmult36} {iopath_Amult1_Cmult37} {iopath_Amult1_Cmult38} {iopath_Amult1_Cmult39} {iopath_Amult1_Cmult40} {iopath_Amult1_Cmult41} {iopath_Amult1_Cmult42} {iopath_Amult1_Cmult43} {iopath_Amult1_Cmult44} {iopath_Amult1_Cmult45} {iopath_Amult1_Cmult46} {iopath_Amult1_Cmult47} {iopath_Amult1_Cmult48} {iopath_Amult1_Cmult49} {iopath_Amult1_Cmult50} {iopath_Amult1_Cmult51} {iopath_Amult1_Cmult52} {iopath_Amult1_Cmult53} {iopath_Amult1_Cmult54} {iopath_Amult1_Cmult55} {iopath_Amult1_Cmult56} {iopath_Amult1_Cmult57} {iopath_Amult1_Cmult58} {iopath_Amult1_Cmult59} {iopath_Amult1_Cmult60} {iopath_Amult1_Cmult61} {iopath_Amult1_Cmult62} {iopath_Amult1_Cmult63} 0 0 {iopath_Amult2_Cmult2} {iopath_Amult2_Cmult3} {iopath_Amult2_Cmult4} {iopath_Amult2_Cmult5} {iopath_Amult2_Cmult6} {iopath_Amult2_Cmult7} {iopath_Amult2_Cmult8} {iopath_Amult2_Cmult9} {iopath_Amult2_Cmult10} {iopath_Amult2_Cmult11} {iopath_Amult2_Cmult12} {iopath_Amult2_Cmult13} {iopath_Amult2_Cmult14} {iopath_Amult2_Cmult15} {iopath_Amult2_Cmult16} {iopath_Amult2_Cmult17} {iopath_Amult2_Cmult18} {iopath_Amult2_Cmult19} {iopath_Amult2_Cmult20} {iopath_Amult2_Cmult21} {iopath_Amult2_Cmult22} {iopath_Amult2_Cmult23} {iopath_Amult2_Cmult24} {iopath_Amult2_Cmult25} {iopath_Amult2_Cmult26} {iopath_Amult2_Cmult27} {iopath_Amult2_Cmult28} {iopath_Amult2_Cmult29} {iopath_Amult2_Cmult30} {iopath_Amult2_Cmult31} {iopath_Amult2_Cmult32} {iopath_Amult2_Cmult33} {iopath_Amult2_Cmult34} {iopath_Amult2_Cmult35} {iopath_Amult2_Cmult36} {iopath_Amult2_Cmult37} {iopath_Amult2_Cmult38} {iopath_Amult2_Cmult39} {iopath_Amult2_Cmult40} {iopath_Amult2_Cmult41} {iopath_Amult2_Cmult42} {iopath_Amult2_Cmult43} {iopath_Amult2_Cmult44} {iopath_Amult2_Cmult45} {iopath_Amult2_Cmult46} {iopath_Amult2_Cmult47} {iopath_Amult2_Cmult48} {iopath_Amult2_Cmult49} {iopath_Amult2_Cmult50} {iopath_Amult2_Cmult51} {iopath_Amult2_Cmult52} {iopath_Amult2_Cmult53} {iopath_Amult2_Cmult54} {iopath_Amult2_Cmult55} {iopath_Amult2_Cmult56} {iopath_Amult2_Cmult57} {iopath_Amult2_Cmult58} {iopath_Amult2_Cmult59} {iopath_Amult2_Cmult60} {iopath_Amult2_Cmult61} {iopath_Amult2_Cmult62} {iopath_Amult2_Cmult63} 0 0 0 {iopath_Amult3_Cmult3} {iopath_Amult3_Cmult4} {iopath_Amult3_Cmult5} {iopath_Amult3_Cmult6} {iopath_Amult3_Cmult7} {iopath_Amult3_Cmult8} {iopath_Amult3_Cmult9} {iopath_Amult3_Cmult10} {iopath_Amult3_Cmult11} {iopath_Amult3_Cmult12} {iopath_Amult3_Cmult13} {iopath_Amult3_Cmult14} {iopath_Amult3_Cmult15} {iopath_Amult3_Cmult16} {iopath_Amult3_Cmult17} {iopath_Amult3_Cmult18} {iopath_Amult3_Cmult19} {iopath_Amult3_Cmult20} {iopath_Amult3_Cmult21} {iopath_Amult3_Cmult22} {iopath_Amult3_Cmult23} {iopath_Amult3_Cmult24} {iopath_Amult3_Cmult25} {iopath_Amult3_Cmult26} {iopath_Amult3_Cmult27} {iopath_Amult3_Cmult28} {iopath_Amult3_Cmult29} {iopath_Amult3_Cmult30} {iopath_Amult3_Cmult31} {iopath_Amult3_Cmult32} {iopath_Amult3_Cmult33} {iopath_Amult3_Cmult34} {iopath_Amult3_Cmult35} {iopath_Amult3_Cmult36} {iopath_Amult3_Cmult37} {iopath_Amult3_Cmult38} {iopath_Amult3_Cmult39} {iopath_Amult3_Cmult40} {iopath_Amult3_Cmult41} {iopath_Amult3_Cmult42} {iopath_Amult3_Cmult43} {iopath_Amult3_Cmult44} {iopath_Amult3_Cmult45} {iopath_Amult3_Cmult46} {iopath_Amult3_Cmult47} {iopath_Amult3_Cmult48} {iopath_Amult3_Cmult49} {iopath_Amult3_Cmult50} {iopath_Amult3_Cmult51} {iopath_Amult3_Cmult52} {iopath_Amult3_Cmult53} {iopath_Amult3_Cmult54} {iopath_Amult3_Cmult55} {iopath_Amult3_Cmult56} {iopath_Amult3_Cmult57} {iopath_Amult3_Cmult58} {iopath_Amult3_Cmult59} {iopath_Amult3_Cmult60} {iopath_Amult3_Cmult61} {iopath_Amult3_Cmult62} {iopath_Amult3_Cmult63} 0 0 0 0 {iopath_Amult4_Cmult4} {iopath_Amult4_Cmult5} {iopath_Amult4_Cmult6} {iopath_Amult4_Cmult7} {iopath_Amult4_Cmult8} {iopath_Amult4_Cmult9} {iopath_Amult4_Cmult10} {iopath_Amult4_Cmult11} {iopath_Amult4_Cmult12} {iopath_Amult4_Cmult13} {iopath_Amult4_Cmult14} {iopath_Amult4_Cmult15} {iopath_Amult4_Cmult16} {iopath_Amult4_Cmult17} {iopath_Amult4_Cmult18} {iopath_Amult4_Cmult19} {iopath_Amult4_Cmult20} {iopath_Amult4_Cmult21} {iopath_Amult4_Cmult22} {iopath_Amult4_Cmult23} {iopath_Amult4_Cmult24} {iopath_Amult4_Cmult25} {iopath_Amult4_Cmult26} {iopath_Amult4_Cmult27} {iopath_Amult4_Cmult28} {iopath_Amult4_Cmult29} {iopath_Amult4_Cmult30} {iopath_Amult4_Cmult31} {iopath_Amult4_Cmult32} {iopath_Amult4_Cmult33} {iopath_Amult4_Cmult34} {iopath_Amult4_Cmult35} {iopath_Amult4_Cmult36} {iopath_Amult4_Cmult37} {iopath_Amult4_Cmult38} {iopath_Amult4_Cmult39} {iopath_Amult4_Cmult40} {iopath_Amult4_Cmult41} {iopath_Amult4_Cmult42} {iopath_Amult4_Cmult43} {iopath_Amult4_Cmult44} {iopath_Amult4_Cmult45} {iopath_Amult4_Cmult46} {iopath_Amult4_Cmult47} {iopath_Amult4_Cmult48} {iopath_Amult4_Cmult49} {iopath_Amult4_Cmult50} {iopath_Amult4_Cmult51} {iopath_Amult4_Cmult52} {iopath_Amult4_Cmult53} {iopath_Amult4_Cmult54} {iopath_Amult4_Cmult55} {iopath_Amult4_Cmult56} {iopath_Amult4_Cmult57} {iopath_Amult4_Cmult58} {iopath_Amult4_Cmult59} {iopath_Amult4_Cmult60} {iopath_Amult4_Cmult61} {iopath_Amult4_Cmult62} {iopath_Amult4_Cmult63} 0 0 0 0 0 {iopath_Amult5_Cmult5} {iopath_Amult5_Cmult6} {iopath_Amult5_Cmult7} {iopath_Amult5_Cmult8} {iopath_Amult5_Cmult9} {iopath_Amult5_Cmult10} {iopath_Amult5_Cmult11} {iopath_Amult5_Cmult12} {iopath_Amult5_Cmult13} {iopath_Amult5_Cmult14} {iopath_Amult5_Cmult15} {iopath_Amult5_Cmult16} {iopath_Amult5_Cmult17} {iopath_Amult5_Cmult18} {iopath_Amult5_Cmult19} {iopath_Amult5_Cmult20} {iopath_Amult5_Cmult21} {iopath_Amult5_Cmult22} {iopath_Amult5_Cmult23} {iopath_Amult5_Cmult24} {iopath_Amult5_Cmult25} {iopath_Amult5_Cmult26} {iopath_Amult5_Cmult27} {iopath_Amult5_Cmult28} {iopath_Amult5_Cmult29} {iopath_Amult5_Cmult30} {iopath_Amult5_Cmult31} {iopath_Amult5_Cmult32} {iopath_Amult5_Cmult33} {iopath_Amult5_Cmult34} {iopath_Amult5_Cmult35} {iopath_Amult5_Cmult36} {iopath_Amult5_Cmult37} {iopath_Amult5_Cmult38} {iopath_Amult5_Cmult39} {iopath_Amult5_Cmult40} {iopath_Amult5_Cmult41} {iopath_Amult5_Cmult42} {iopath_Amult5_Cmult43} {iopath_Amult5_Cmult44} {iopath_Amult5_Cmult45} {iopath_Amult5_Cmult46} {iopath_Amult5_Cmult47} {iopath_Amult5_Cmult48} {iopath_Amult5_Cmult49} {iopath_Amult5_Cmult50} {iopath_Amult5_Cmult51} {iopath_Amult5_Cmult52} {iopath_Amult5_Cmult53} {iopath_Amult5_Cmult54} {iopath_Amult5_Cmult55} {iopath_Amult5_Cmult56} {iopath_Amult5_Cmult57} {iopath_Amult5_Cmult58} {iopath_Amult5_Cmult59} {iopath_Amult5_Cmult60} {iopath_Amult5_Cmult61} {iopath_Amult5_Cmult62} {iopath_Amult5_Cmult63} 0 0 0 0 0 0 {iopath_Amult6_Cmult6} {iopath_Amult6_Cmult7} {iopath_Amult6_Cmult8} {iopath_Amult6_Cmult9} {iopath_Amult6_Cmult10} {iopath_Amult6_Cmult11} {iopath_Amult6_Cmult12} {iopath_Amult6_Cmult13} {iopath_Amult6_Cmult14} {iopath_Amult6_Cmult15} {iopath_Amult6_Cmult16} {iopath_Amult6_Cmult17} {iopath_Amult6_Cmult18} {iopath_Amult6_Cmult19} {iopath_Amult6_Cmult20} {iopath_Amult6_Cmult21} {iopath_Amult6_Cmult22} {iopath_Amult6_Cmult23} {iopath_Amult6_Cmult24} {iopath_Amult6_Cmult25} {iopath_Amult6_Cmult26} {iopath_Amult6_Cmult27} {iopath_Amult6_Cmult28} {iopath_Amult6_Cmult29} {iopath_Amult6_Cmult30} {iopath_Amult6_Cmult31} {iopath_Amult6_Cmult32} {iopath_Amult6_Cmult33} {iopath_Amult6_Cmult34} {iopath_Amult6_Cmult35} {iopath_Amult6_Cmult36} {iopath_Amult6_Cmult37} {iopath_Amult6_Cmult38} {iopath_Amult6_Cmult39} {iopath_Amult6_Cmult40} {iopath_Amult6_Cmult41} {iopath_Amult6_Cmult42} {iopath_Amult6_Cmult43} {iopath_Amult6_Cmult44} {iopath_Amult6_Cmult45} {iopath_Amult6_Cmult46} {iopath_Amult6_Cmult47} {iopath_Amult6_Cmult48} {iopath_Amult6_Cmult49} {iopath_Amult6_Cmult50} {iopath_Amult6_Cmult51} {iopath_Amult6_Cmult52} {iopath_Amult6_Cmult53} {iopath_Amult6_Cmult54} {iopath_Amult6_Cmult55} {iopath_Amult6_Cmult56} {iopath_Amult6_Cmult57} {iopath_Amult6_Cmult58} {iopath_Amult6_Cmult59} {iopath_Amult6_Cmult60} {iopath_Amult6_Cmult61} {iopath_Amult6_Cmult62} {iopath_Amult6_Cmult63} 0 0 0 0 0 0 0 {iopath_Amult7_Cmult7} {iopath_Amult7_Cmult8} {iopath_Amult7_Cmult9} {iopath_Amult7_Cmult10} {iopath_Amult7_Cmult11} {iopath_Amult7_Cmult12} {iopath_Amult7_Cmult13} {iopath_Amult7_Cmult14} {iopath_Amult7_Cmult15} {iopath_Amult7_Cmult16} {iopath_Amult7_Cmult17} {iopath_Amult7_Cmult18} {iopath_Amult7_Cmult19} {iopath_Amult7_Cmult20} {iopath_Amult7_Cmult21} {iopath_Amult7_Cmult22} {iopath_Amult7_Cmult23} {iopath_Amult7_Cmult24} {iopath_Amult7_Cmult25} {iopath_Amult7_Cmult26} {iopath_Amult7_Cmult27} {iopath_Amult7_Cmult28} {iopath_Amult7_Cmult29} {iopath_Amult7_Cmult30} {iopath_Amult7_Cmult31} {iopath_Amult7_Cmult32} {iopath_Amult7_Cmult33} {iopath_Amult7_Cmult34} {iopath_Amult7_Cmult35} {iopath_Amult7_Cmult36} {iopath_Amult7_Cmult37} {iopath_Amult7_Cmult38} {iopath_Amult7_Cmult39} {iopath_Amult7_Cmult40} {iopath_Amult7_Cmult41} {iopath_Amult7_Cmult42} {iopath_Amult7_Cmult43} {iopath_Amult7_Cmult44} {iopath_Amult7_Cmult45} {iopath_Amult7_Cmult46} {iopath_Amult7_Cmult47} {iopath_Amult7_Cmult48} {iopath_Amult7_Cmult49} {iopath_Amult7_Cmult50} {iopath_Amult7_Cmult51} {iopath_Amult7_Cmult52} {iopath_Amult7_Cmult53} {iopath_Amult7_Cmult54} {iopath_Amult7_Cmult55} {iopath_Amult7_Cmult56} {iopath_Amult7_Cmult57} {iopath_Amult7_Cmult58} {iopath_Amult7_Cmult59} {iopath_Amult7_Cmult60} {iopath_Amult7_Cmult61} {iopath_Amult7_Cmult62} {iopath_Amult7_Cmult63} 0 0 0 0 0 0 0 0 {iopath_Amult8_Cmult8} {iopath_Amult8_Cmult9} {iopath_Amult8_Cmult10} {iopath_Amult8_Cmult11} {iopath_Amult8_Cmult12} {iopath_Amult8_Cmult13} {iopath_Amult8_Cmult14} {iopath_Amult8_Cmult15} {iopath_Amult8_Cmult16} {iopath_Amult8_Cmult17} {iopath_Amult8_Cmult18} {iopath_Amult8_Cmult19} {iopath_Amult8_Cmult20} {iopath_Amult8_Cmult21} {iopath_Amult8_Cmult22} {iopath_Amult8_Cmult23} {iopath_Amult8_Cmult24} {iopath_Amult8_Cmult25} {iopath_Amult8_Cmult26} {iopath_Amult8_Cmult27} {iopath_Amult8_Cmult28} {iopath_Amult8_Cmult29} {iopath_Amult8_Cmult30} {iopath_Amult8_Cmult31} {iopath_Amult8_Cmult32} {iopath_Amult8_Cmult33} {iopath_Amult8_Cmult34} {iopath_Amult8_Cmult35} {iopath_Amult8_Cmult36} {iopath_Amult8_Cmult37} {iopath_Amult8_Cmult38} {iopath_Amult8_Cmult39} {iopath_Amult8_Cmult40} {iopath_Amult8_Cmult41} {iopath_Amult8_Cmult42} {iopath_Amult8_Cmult43} {iopath_Amult8_Cmult44} {iopath_Amult8_Cmult45} {iopath_Amult8_Cmult46} {iopath_Amult8_Cmult47} {iopath_Amult8_Cmult48} {iopath_Amult8_Cmult49} {iopath_Amult8_Cmult50} {iopath_Amult8_Cmult51} {iopath_Amult8_Cmult52} {iopath_Amult8_Cmult53} {iopath_Amult8_Cmult54} {iopath_Amult8_Cmult55} {iopath_Amult8_Cmult56} {iopath_Amult8_Cmult57} {iopath_Amult8_Cmult58} {iopath_Amult8_Cmult59} {iopath_Amult8_Cmult60} {iopath_Amult8_Cmult61} {iopath_Amult8_Cmult62} {iopath_Amult8_Cmult63} 0 0 0 0 0 0 0 0 0 {iopath_Amult9_Cmult9} {iopath_Amult9_Cmult10} {iopath_Amult9_Cmult11} {iopath_Amult9_Cmult12} {iopath_Amult9_Cmult13} {iopath_Amult9_Cmult14} {iopath_Amult9_Cmult15} {iopath_Amult9_Cmult16} {iopath_Amult9_Cmult17} {iopath_Amult9_Cmult18} {iopath_Amult9_Cmult19} {iopath_Amult9_Cmult20} {iopath_Amult9_Cmult21} {iopath_Amult9_Cmult22} {iopath_Amult9_Cmult23} {iopath_Amult9_Cmult24} {iopath_Amult9_Cmult25} {iopath_Amult9_Cmult26} {iopath_Amult9_Cmult27} {iopath_Amult9_Cmult28} {iopath_Amult9_Cmult29} {iopath_Amult9_Cmult30} {iopath_Amult9_Cmult31} {iopath_Amult9_Cmult32} {iopath_Amult9_Cmult33} {iopath_Amult9_Cmult34} {iopath_Amult9_Cmult35} {iopath_Amult9_Cmult36} {iopath_Amult9_Cmult37} {iopath_Amult9_Cmult38} {iopath_Amult9_Cmult39} {iopath_Amult9_Cmult40} {iopath_Amult9_Cmult41} {iopath_Amult9_Cmult42} {iopath_Amult9_Cmult43} {iopath_Amult9_Cmult44} {iopath_Amult9_Cmult45} {iopath_Amult9_Cmult46} {iopath_Amult9_Cmult47} {iopath_Amult9_Cmult48} {iopath_Amult9_Cmult49} {iopath_Amult9_Cmult50} {iopath_Amult9_Cmult51} {iopath_Amult9_Cmult52} {iopath_Amult9_Cmult53} {iopath_Amult9_Cmult54} {iopath_Amult9_Cmult55} {iopath_Amult9_Cmult56} {iopath_Amult9_Cmult57} {iopath_Amult9_Cmult58} {iopath_Amult9_Cmult59} {iopath_Amult9_Cmult60} {iopath_Amult9_Cmult61} {iopath_Amult9_Cmult62} {iopath_Amult9_Cmult63} 0 0 0 0 0 0 0 0 0 0 {iopath_Amult10_Cmult10} {iopath_Amult10_Cmult11} {iopath_Amult10_Cmult12} {iopath_Amult10_Cmult13} {iopath_Amult10_Cmult14} {iopath_Amult10_Cmult15} {iopath_Amult10_Cmult16} {iopath_Amult10_Cmult17} {iopath_Amult10_Cmult18} {iopath_Amult10_Cmult19} {iopath_Amult10_Cmult20} {iopath_Amult10_Cmult21} {iopath_Amult10_Cmult22} {iopath_Amult10_Cmult23} {iopath_Amult10_Cmult24} {iopath_Amult10_Cmult25} {iopath_Amult10_Cmult26} {iopath_Amult10_Cmult27} {iopath_Amult10_Cmult28} {iopath_Amult10_Cmult29} {iopath_Amult10_Cmult30} {iopath_Amult10_Cmult31} {iopath_Amult10_Cmult32} {iopath_Amult10_Cmult33} {iopath_Amult10_Cmult34} {iopath_Amult10_Cmult35} {iopath_Amult10_Cmult36} {iopath_Amult10_Cmult37} {iopath_Amult10_Cmult38} {iopath_Amult10_Cmult39} {iopath_Amult10_Cmult40} {iopath_Amult10_Cmult41} {iopath_Amult10_Cmult42} {iopath_Amult10_Cmult43} {iopath_Amult10_Cmult44} {iopath_Amult10_Cmult45} {iopath_Amult10_Cmult46} {iopath_Amult10_Cmult47} {iopath_Amult10_Cmult48} {iopath_Amult10_Cmult49} {iopath_Amult10_Cmult50} {iopath_Amult10_Cmult51} {iopath_Amult10_Cmult52} {iopath_Amult10_Cmult53} {iopath_Amult10_Cmult54} {iopath_Amult10_Cmult55} {iopath_Amult10_Cmult56} {iopath_Amult10_Cmult57} {iopath_Amult10_Cmult58} {iopath_Amult10_Cmult59} {iopath_Amult10_Cmult60} {iopath_Amult10_Cmult61} {iopath_Amult10_Cmult62} {iopath_Amult10_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult11_Cmult11} {iopath_Amult11_Cmult12} {iopath_Amult11_Cmult13} {iopath_Amult11_Cmult14} {iopath_Amult11_Cmult15} {iopath_Amult11_Cmult16} {iopath_Amult11_Cmult17} {iopath_Amult11_Cmult18} {iopath_Amult11_Cmult19} {iopath_Amult11_Cmult20} {iopath_Amult11_Cmult21} {iopath_Amult11_Cmult22} {iopath_Amult11_Cmult23} {iopath_Amult11_Cmult24} {iopath_Amult11_Cmult25} {iopath_Amult11_Cmult26} {iopath_Amult11_Cmult27} {iopath_Amult11_Cmult28} {iopath_Amult11_Cmult29} {iopath_Amult11_Cmult30} {iopath_Amult11_Cmult31} {iopath_Amult11_Cmult32} {iopath_Amult11_Cmult33} {iopath_Amult11_Cmult34} {iopath_Amult11_Cmult35} {iopath_Amult11_Cmult36} {iopath_Amult11_Cmult37} {iopath_Amult11_Cmult38} {iopath_Amult11_Cmult39} {iopath_Amult11_Cmult40} {iopath_Amult11_Cmult41} {iopath_Amult11_Cmult42} {iopath_Amult11_Cmult43} {iopath_Amult11_Cmult44} {iopath_Amult11_Cmult45} {iopath_Amult11_Cmult46} {iopath_Amult11_Cmult47} {iopath_Amult11_Cmult48} {iopath_Amult11_Cmult49} {iopath_Amult11_Cmult50} {iopath_Amult11_Cmult51} {iopath_Amult11_Cmult52} {iopath_Amult11_Cmult53} {iopath_Amult11_Cmult54} {iopath_Amult11_Cmult55} {iopath_Amult11_Cmult56} {iopath_Amult11_Cmult57} {iopath_Amult11_Cmult58} {iopath_Amult11_Cmult59} {iopath_Amult11_Cmult60} {iopath_Amult11_Cmult61} {iopath_Amult11_Cmult62} {iopath_Amult11_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult12_Cmult12} {iopath_Amult12_Cmult13} {iopath_Amult12_Cmult14} {iopath_Amult12_Cmult15} {iopath_Amult12_Cmult16} {iopath_Amult12_Cmult17} {iopath_Amult12_Cmult18} {iopath_Amult12_Cmult19} {iopath_Amult12_Cmult20} {iopath_Amult12_Cmult21} {iopath_Amult12_Cmult22} {iopath_Amult12_Cmult23} {iopath_Amult12_Cmult24} {iopath_Amult12_Cmult25} {iopath_Amult12_Cmult26} {iopath_Amult12_Cmult27} {iopath_Amult12_Cmult28} {iopath_Amult12_Cmult29} {iopath_Amult12_Cmult30} {iopath_Amult12_Cmult31} {iopath_Amult12_Cmult32} {iopath_Amult12_Cmult33} {iopath_Amult12_Cmult34} {iopath_Amult12_Cmult35} {iopath_Amult12_Cmult36} {iopath_Amult12_Cmult37} {iopath_Amult12_Cmult38} {iopath_Amult12_Cmult39} {iopath_Amult12_Cmult40} {iopath_Amult12_Cmult41} {iopath_Amult12_Cmult42} {iopath_Amult12_Cmult43} {iopath_Amult12_Cmult44} {iopath_Amult12_Cmult45} {iopath_Amult12_Cmult46} {iopath_Amult12_Cmult47} {iopath_Amult12_Cmult48} {iopath_Amult12_Cmult49} {iopath_Amult12_Cmult50} {iopath_Amult12_Cmult51} {iopath_Amult12_Cmult52} {iopath_Amult12_Cmult53} {iopath_Amult12_Cmult54} {iopath_Amult12_Cmult55} {iopath_Amult12_Cmult56} {iopath_Amult12_Cmult57} {iopath_Amult12_Cmult58} {iopath_Amult12_Cmult59} {iopath_Amult12_Cmult60} {iopath_Amult12_Cmult61} {iopath_Amult12_Cmult62} {iopath_Amult12_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult13_Cmult13} {iopath_Amult13_Cmult14} {iopath_Amult13_Cmult15} {iopath_Amult13_Cmult16} {iopath_Amult13_Cmult17} {iopath_Amult13_Cmult18} {iopath_Amult13_Cmult19} {iopath_Amult13_Cmult20} {iopath_Amult13_Cmult21} {iopath_Amult13_Cmult22} {iopath_Amult13_Cmult23} {iopath_Amult13_Cmult24} {iopath_Amult13_Cmult25} {iopath_Amult13_Cmult26} {iopath_Amult13_Cmult27} {iopath_Amult13_Cmult28} {iopath_Amult13_Cmult29} {iopath_Amult13_Cmult30} {iopath_Amult13_Cmult31} {iopath_Amult13_Cmult32} {iopath_Amult13_Cmult33} {iopath_Amult13_Cmult34} {iopath_Amult13_Cmult35} {iopath_Amult13_Cmult36} {iopath_Amult13_Cmult37} {iopath_Amult13_Cmult38} {iopath_Amult13_Cmult39} {iopath_Amult13_Cmult40} {iopath_Amult13_Cmult41} {iopath_Amult13_Cmult42} {iopath_Amult13_Cmult43} {iopath_Amult13_Cmult44} {iopath_Amult13_Cmult45} {iopath_Amult13_Cmult46} {iopath_Amult13_Cmult47} {iopath_Amult13_Cmult48} {iopath_Amult13_Cmult49} {iopath_Amult13_Cmult50} {iopath_Amult13_Cmult51} {iopath_Amult13_Cmult52} {iopath_Amult13_Cmult53} {iopath_Amult13_Cmult54} {iopath_Amult13_Cmult55} {iopath_Amult13_Cmult56} {iopath_Amult13_Cmult57} {iopath_Amult13_Cmult58} {iopath_Amult13_Cmult59} {iopath_Amult13_Cmult60} {iopath_Amult13_Cmult61} {iopath_Amult13_Cmult62} {iopath_Amult13_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult14_Cmult14} {iopath_Amult14_Cmult15} {iopath_Amult14_Cmult16} {iopath_Amult14_Cmult17} {iopath_Amult14_Cmult18} {iopath_Amult14_Cmult19} {iopath_Amult14_Cmult20} {iopath_Amult14_Cmult21} {iopath_Amult14_Cmult22} {iopath_Amult14_Cmult23} {iopath_Amult14_Cmult24} {iopath_Amult14_Cmult25} {iopath_Amult14_Cmult26} {iopath_Amult14_Cmult27} {iopath_Amult14_Cmult28} {iopath_Amult14_Cmult29} {iopath_Amult14_Cmult30} {iopath_Amult14_Cmult31} {iopath_Amult14_Cmult32} {iopath_Amult14_Cmult33} {iopath_Amult14_Cmult34} {iopath_Amult14_Cmult35} {iopath_Amult14_Cmult36} {iopath_Amult14_Cmult37} {iopath_Amult14_Cmult38} {iopath_Amult14_Cmult39} {iopath_Amult14_Cmult40} {iopath_Amult14_Cmult41} {iopath_Amult14_Cmult42} {iopath_Amult14_Cmult43} {iopath_Amult14_Cmult44} {iopath_Amult14_Cmult45} {iopath_Amult14_Cmult46} {iopath_Amult14_Cmult47} {iopath_Amult14_Cmult48} {iopath_Amult14_Cmult49} {iopath_Amult14_Cmult50} {iopath_Amult14_Cmult51} {iopath_Amult14_Cmult52} {iopath_Amult14_Cmult53} {iopath_Amult14_Cmult54} {iopath_Amult14_Cmult55} {iopath_Amult14_Cmult56} {iopath_Amult14_Cmult57} {iopath_Amult14_Cmult58} {iopath_Amult14_Cmult59} {iopath_Amult14_Cmult60} {iopath_Amult14_Cmult61} {iopath_Amult14_Cmult62} {iopath_Amult14_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult15_Cmult15} {iopath_Amult15_Cmult16} {iopath_Amult15_Cmult17} {iopath_Amult15_Cmult18} {iopath_Amult15_Cmult19} {iopath_Amult15_Cmult20} {iopath_Amult15_Cmult21} {iopath_Amult15_Cmult22} {iopath_Amult15_Cmult23} {iopath_Amult15_Cmult24} {iopath_Amult15_Cmult25} {iopath_Amult15_Cmult26} {iopath_Amult15_Cmult27} {iopath_Amult15_Cmult28} {iopath_Amult15_Cmult29} {iopath_Amult15_Cmult30} {iopath_Amult15_Cmult31} {iopath_Amult15_Cmult32} {iopath_Amult15_Cmult33} {iopath_Amult15_Cmult34} {iopath_Amult15_Cmult35} {iopath_Amult15_Cmult36} {iopath_Amult15_Cmult37} {iopath_Amult15_Cmult38} {iopath_Amult15_Cmult39} {iopath_Amult15_Cmult40} {iopath_Amult15_Cmult41} {iopath_Amult15_Cmult42} {iopath_Amult15_Cmult43} {iopath_Amult15_Cmult44} {iopath_Amult15_Cmult45} {iopath_Amult15_Cmult46} {iopath_Amult15_Cmult47} {iopath_Amult15_Cmult48} {iopath_Amult15_Cmult49} {iopath_Amult15_Cmult50} {iopath_Amult15_Cmult51} {iopath_Amult15_Cmult52} {iopath_Amult15_Cmult53} {iopath_Amult15_Cmult54} {iopath_Amult15_Cmult55} {iopath_Amult15_Cmult56} {iopath_Amult15_Cmult57} {iopath_Amult15_Cmult58} {iopath_Amult15_Cmult59} {iopath_Amult15_Cmult60} {iopath_Amult15_Cmult61} {iopath_Amult15_Cmult62} {iopath_Amult15_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult16_Cmult16} {iopath_Amult16_Cmult17} {iopath_Amult16_Cmult18} {iopath_Amult16_Cmult19} {iopath_Amult16_Cmult20} {iopath_Amult16_Cmult21} {iopath_Amult16_Cmult22} {iopath_Amult16_Cmult23} {iopath_Amult16_Cmult24} {iopath_Amult16_Cmult25} {iopath_Amult16_Cmult26} {iopath_Amult16_Cmult27} {iopath_Amult16_Cmult28} {iopath_Amult16_Cmult29} {iopath_Amult16_Cmult30} {iopath_Amult16_Cmult31} {iopath_Amult16_Cmult32} {iopath_Amult16_Cmult33} {iopath_Amult16_Cmult34} {iopath_Amult16_Cmult35} {iopath_Amult16_Cmult36} {iopath_Amult16_Cmult37} {iopath_Amult16_Cmult38} {iopath_Amult16_Cmult39} {iopath_Amult16_Cmult40} {iopath_Amult16_Cmult41} {iopath_Amult16_Cmult42} {iopath_Amult16_Cmult43} {iopath_Amult16_Cmult44} {iopath_Amult16_Cmult45} {iopath_Amult16_Cmult46} {iopath_Amult16_Cmult47} {iopath_Amult16_Cmult48} {iopath_Amult16_Cmult49} {iopath_Amult16_Cmult50} {iopath_Amult16_Cmult51} {iopath_Amult16_Cmult52} {iopath_Amult16_Cmult53} {iopath_Amult16_Cmult54} {iopath_Amult16_Cmult55} {iopath_Amult16_Cmult56} {iopath_Amult16_Cmult57} {iopath_Amult16_Cmult58} {iopath_Amult16_Cmult59} {iopath_Amult16_Cmult60} {iopath_Amult16_Cmult61} {iopath_Amult16_Cmult62} {iopath_Amult16_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult17_Cmult17} {iopath_Amult17_Cmult18} {iopath_Amult17_Cmult19} {iopath_Amult17_Cmult20} {iopath_Amult17_Cmult21} {iopath_Amult17_Cmult22} {iopath_Amult17_Cmult23} {iopath_Amult17_Cmult24} {iopath_Amult17_Cmult25} {iopath_Amult17_Cmult26} {iopath_Amult17_Cmult27} {iopath_Amult17_Cmult28} {iopath_Amult17_Cmult29} {iopath_Amult17_Cmult30} {iopath_Amult17_Cmult31} {iopath_Amult17_Cmult32} {iopath_Amult17_Cmult33} {iopath_Amult17_Cmult34} {iopath_Amult17_Cmult35} {iopath_Amult17_Cmult36} {iopath_Amult17_Cmult37} {iopath_Amult17_Cmult38} {iopath_Amult17_Cmult39} {iopath_Amult17_Cmult40} {iopath_Amult17_Cmult41} {iopath_Amult17_Cmult42} {iopath_Amult17_Cmult43} {iopath_Amult17_Cmult44} {iopath_Amult17_Cmult45} {iopath_Amult17_Cmult46} {iopath_Amult17_Cmult47} {iopath_Amult17_Cmult48} {iopath_Amult17_Cmult49} {iopath_Amult17_Cmult50} {iopath_Amult17_Cmult51} {iopath_Amult17_Cmult52} {iopath_Amult17_Cmult53} {iopath_Amult17_Cmult54} {iopath_Amult17_Cmult55} {iopath_Amult17_Cmult56} {iopath_Amult17_Cmult57} {iopath_Amult17_Cmult58} {iopath_Amult17_Cmult59} {iopath_Amult17_Cmult60} {iopath_Amult17_Cmult61} {iopath_Amult17_Cmult62} {iopath_Amult17_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult18_Cmult18} {iopath_Amult18_Cmult19} {iopath_Amult18_Cmult20} {iopath_Amult18_Cmult21} {iopath_Amult18_Cmult22} {iopath_Amult18_Cmult23} {iopath_Amult18_Cmult24} {iopath_Amult18_Cmult25} {iopath_Amult18_Cmult26} {iopath_Amult18_Cmult27} {iopath_Amult18_Cmult28} {iopath_Amult18_Cmult29} {iopath_Amult18_Cmult30} {iopath_Amult18_Cmult31} {iopath_Amult18_Cmult32} {iopath_Amult18_Cmult33} {iopath_Amult18_Cmult34} {iopath_Amult18_Cmult35} {iopath_Amult18_Cmult36} {iopath_Amult18_Cmult37} {iopath_Amult18_Cmult38} {iopath_Amult18_Cmult39} {iopath_Amult18_Cmult40} {iopath_Amult18_Cmult41} {iopath_Amult18_Cmult42} {iopath_Amult18_Cmult43} {iopath_Amult18_Cmult44} {iopath_Amult18_Cmult45} {iopath_Amult18_Cmult46} {iopath_Amult18_Cmult47} {iopath_Amult18_Cmult48} {iopath_Amult18_Cmult49} {iopath_Amult18_Cmult50} {iopath_Amult18_Cmult51} {iopath_Amult18_Cmult52} {iopath_Amult18_Cmult53} {iopath_Amult18_Cmult54} {iopath_Amult18_Cmult55} {iopath_Amult18_Cmult56} {iopath_Amult18_Cmult57} {iopath_Amult18_Cmult58} {iopath_Amult18_Cmult59} {iopath_Amult18_Cmult60} {iopath_Amult18_Cmult61} {iopath_Amult18_Cmult62} {iopath_Amult18_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult19_Cmult19} {iopath_Amult19_Cmult20} {iopath_Amult19_Cmult21} {iopath_Amult19_Cmult22} {iopath_Amult19_Cmult23} {iopath_Amult19_Cmult24} {iopath_Amult19_Cmult25} {iopath_Amult19_Cmult26} {iopath_Amult19_Cmult27} {iopath_Amult19_Cmult28} {iopath_Amult19_Cmult29} {iopath_Amult19_Cmult30} {iopath_Amult19_Cmult31} {iopath_Amult19_Cmult32} {iopath_Amult19_Cmult33} {iopath_Amult19_Cmult34} {iopath_Amult19_Cmult35} {iopath_Amult19_Cmult36} {iopath_Amult19_Cmult37} {iopath_Amult19_Cmult38} {iopath_Amult19_Cmult39} {iopath_Amult19_Cmult40} {iopath_Amult19_Cmult41} {iopath_Amult19_Cmult42} {iopath_Amult19_Cmult43} {iopath_Amult19_Cmult44} {iopath_Amult19_Cmult45} {iopath_Amult19_Cmult46} {iopath_Amult19_Cmult47} {iopath_Amult19_Cmult48} {iopath_Amult19_Cmult49} {iopath_Amult19_Cmult50} {iopath_Amult19_Cmult51} {iopath_Amult19_Cmult52} {iopath_Amult19_Cmult53} {iopath_Amult19_Cmult54} {iopath_Amult19_Cmult55} {iopath_Amult19_Cmult56} {iopath_Amult19_Cmult57} {iopath_Amult19_Cmult58} {iopath_Amult19_Cmult59} {iopath_Amult19_Cmult60} {iopath_Amult19_Cmult61} {iopath_Amult19_Cmult62} {iopath_Amult19_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult20_Cmult20} {iopath_Amult20_Cmult21} {iopath_Amult20_Cmult22} {iopath_Amult20_Cmult23} {iopath_Amult20_Cmult24} {iopath_Amult20_Cmult25} {iopath_Amult20_Cmult26} {iopath_Amult20_Cmult27} {iopath_Amult20_Cmult28} {iopath_Amult20_Cmult29} {iopath_Amult20_Cmult30} {iopath_Amult20_Cmult31} {iopath_Amult20_Cmult32} {iopath_Amult20_Cmult33} {iopath_Amult20_Cmult34} {iopath_Amult20_Cmult35} {iopath_Amult20_Cmult36} {iopath_Amult20_Cmult37} {iopath_Amult20_Cmult38} {iopath_Amult20_Cmult39} {iopath_Amult20_Cmult40} {iopath_Amult20_Cmult41} {iopath_Amult20_Cmult42} {iopath_Amult20_Cmult43} {iopath_Amult20_Cmult44} {iopath_Amult20_Cmult45} {iopath_Amult20_Cmult46} {iopath_Amult20_Cmult47} {iopath_Amult20_Cmult48} {iopath_Amult20_Cmult49} {iopath_Amult20_Cmult50} {iopath_Amult20_Cmult51} {iopath_Amult20_Cmult52} {iopath_Amult20_Cmult53} {iopath_Amult20_Cmult54} {iopath_Amult20_Cmult55} {iopath_Amult20_Cmult56} {iopath_Amult20_Cmult57} {iopath_Amult20_Cmult58} {iopath_Amult20_Cmult59} {iopath_Amult20_Cmult60} {iopath_Amult20_Cmult61} {iopath_Amult20_Cmult62} {iopath_Amult20_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult21_Cmult21} {iopath_Amult21_Cmult22} {iopath_Amult21_Cmult23} {iopath_Amult21_Cmult24} {iopath_Amult21_Cmult25} {iopath_Amult21_Cmult26} {iopath_Amult21_Cmult27} {iopath_Amult21_Cmult28} {iopath_Amult21_Cmult29} {iopath_Amult21_Cmult30} {iopath_Amult21_Cmult31} {iopath_Amult21_Cmult32} {iopath_Amult21_Cmult33} {iopath_Amult21_Cmult34} {iopath_Amult21_Cmult35} {iopath_Amult21_Cmult36} {iopath_Amult21_Cmult37} {iopath_Amult21_Cmult38} {iopath_Amult21_Cmult39} {iopath_Amult21_Cmult40} {iopath_Amult21_Cmult41} {iopath_Amult21_Cmult42} {iopath_Amult21_Cmult43} {iopath_Amult21_Cmult44} {iopath_Amult21_Cmult45} {iopath_Amult21_Cmult46} {iopath_Amult21_Cmult47} {iopath_Amult21_Cmult48} {iopath_Amult21_Cmult49} {iopath_Amult21_Cmult50} {iopath_Amult21_Cmult51} {iopath_Amult21_Cmult52} {iopath_Amult21_Cmult53} {iopath_Amult21_Cmult54} {iopath_Amult21_Cmult55} {iopath_Amult21_Cmult56} {iopath_Amult21_Cmult57} {iopath_Amult21_Cmult58} {iopath_Amult21_Cmult59} {iopath_Amult21_Cmult60} {iopath_Amult21_Cmult61} {iopath_Amult21_Cmult62} {iopath_Amult21_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult22_Cmult22} {iopath_Amult22_Cmult23} {iopath_Amult22_Cmult24} {iopath_Amult22_Cmult25} {iopath_Amult22_Cmult26} {iopath_Amult22_Cmult27} {iopath_Amult22_Cmult28} {iopath_Amult22_Cmult29} {iopath_Amult22_Cmult30} {iopath_Amult22_Cmult31} {iopath_Amult22_Cmult32} {iopath_Amult22_Cmult33} {iopath_Amult22_Cmult34} {iopath_Amult22_Cmult35} {iopath_Amult22_Cmult36} {iopath_Amult22_Cmult37} {iopath_Amult22_Cmult38} {iopath_Amult22_Cmult39} {iopath_Amult22_Cmult40} {iopath_Amult22_Cmult41} {iopath_Amult22_Cmult42} {iopath_Amult22_Cmult43} {iopath_Amult22_Cmult44} {iopath_Amult22_Cmult45} {iopath_Amult22_Cmult46} {iopath_Amult22_Cmult47} {iopath_Amult22_Cmult48} {iopath_Amult22_Cmult49} {iopath_Amult22_Cmult50} {iopath_Amult22_Cmult51} {iopath_Amult22_Cmult52} {iopath_Amult22_Cmult53} {iopath_Amult22_Cmult54} {iopath_Amult22_Cmult55} {iopath_Amult22_Cmult56} {iopath_Amult22_Cmult57} {iopath_Amult22_Cmult58} {iopath_Amult22_Cmult59} {iopath_Amult22_Cmult60} {iopath_Amult22_Cmult61} {iopath_Amult22_Cmult62} {iopath_Amult22_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult23_Cmult23} {iopath_Amult23_Cmult24} {iopath_Amult23_Cmult25} {iopath_Amult23_Cmult26} {iopath_Amult23_Cmult27} {iopath_Amult23_Cmult28} {iopath_Amult23_Cmult29} {iopath_Amult23_Cmult30} {iopath_Amult23_Cmult31} {iopath_Amult23_Cmult32} {iopath_Amult23_Cmult33} {iopath_Amult23_Cmult34} {iopath_Amult23_Cmult35} {iopath_Amult23_Cmult36} {iopath_Amult23_Cmult37} {iopath_Amult23_Cmult38} {iopath_Amult23_Cmult39} {iopath_Amult23_Cmult40} {iopath_Amult23_Cmult41} {iopath_Amult23_Cmult42} {iopath_Amult23_Cmult43} {iopath_Amult23_Cmult44} {iopath_Amult23_Cmult45} {iopath_Amult23_Cmult46} {iopath_Amult23_Cmult47} {iopath_Amult23_Cmult48} {iopath_Amult23_Cmult49} {iopath_Amult23_Cmult50} {iopath_Amult23_Cmult51} {iopath_Amult23_Cmult52} {iopath_Amult23_Cmult53} {iopath_Amult23_Cmult54} {iopath_Amult23_Cmult55} {iopath_Amult23_Cmult56} {iopath_Amult23_Cmult57} {iopath_Amult23_Cmult58} {iopath_Amult23_Cmult59} {iopath_Amult23_Cmult60} {iopath_Amult23_Cmult61} {iopath_Amult23_Cmult62} {iopath_Amult23_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult24_Cmult24} {iopath_Amult24_Cmult25} {iopath_Amult24_Cmult26} {iopath_Amult24_Cmult27} {iopath_Amult24_Cmult28} {iopath_Amult24_Cmult29} {iopath_Amult24_Cmult30} {iopath_Amult24_Cmult31} {iopath_Amult24_Cmult32} {iopath_Amult24_Cmult33} {iopath_Amult24_Cmult34} {iopath_Amult24_Cmult35} {iopath_Amult24_Cmult36} {iopath_Amult24_Cmult37} {iopath_Amult24_Cmult38} {iopath_Amult24_Cmult39} {iopath_Amult24_Cmult40} {iopath_Amult24_Cmult41} {iopath_Amult24_Cmult42} {iopath_Amult24_Cmult43} {iopath_Amult24_Cmult44} {iopath_Amult24_Cmult45} {iopath_Amult24_Cmult46} {iopath_Amult24_Cmult47} {iopath_Amult24_Cmult48} {iopath_Amult24_Cmult49} {iopath_Amult24_Cmult50} {iopath_Amult24_Cmult51} {iopath_Amult24_Cmult52} {iopath_Amult24_Cmult53} {iopath_Amult24_Cmult54} {iopath_Amult24_Cmult55} {iopath_Amult24_Cmult56} {iopath_Amult24_Cmult57} {iopath_Amult24_Cmult58} {iopath_Amult24_Cmult59} {iopath_Amult24_Cmult60} {iopath_Amult24_Cmult61} {iopath_Amult24_Cmult62} {iopath_Amult24_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult25_Cmult25} {iopath_Amult25_Cmult26} {iopath_Amult25_Cmult27} {iopath_Amult25_Cmult28} {iopath_Amult25_Cmult29} {iopath_Amult25_Cmult30} {iopath_Amult25_Cmult31} {iopath_Amult25_Cmult32} {iopath_Amult25_Cmult33} {iopath_Amult25_Cmult34} {iopath_Amult25_Cmult35} {iopath_Amult25_Cmult36} {iopath_Amult25_Cmult37} {iopath_Amult25_Cmult38} {iopath_Amult25_Cmult39} {iopath_Amult25_Cmult40} {iopath_Amult25_Cmult41} {iopath_Amult25_Cmult42} {iopath_Amult25_Cmult43} {iopath_Amult25_Cmult44} {iopath_Amult25_Cmult45} {iopath_Amult25_Cmult46} {iopath_Amult25_Cmult47} {iopath_Amult25_Cmult48} {iopath_Amult25_Cmult49} {iopath_Amult25_Cmult50} {iopath_Amult25_Cmult51} {iopath_Amult25_Cmult52} {iopath_Amult25_Cmult53} {iopath_Amult25_Cmult54} {iopath_Amult25_Cmult55} {iopath_Amult25_Cmult56} {iopath_Amult25_Cmult57} {iopath_Amult25_Cmult58} {iopath_Amult25_Cmult59} {iopath_Amult25_Cmult60} {iopath_Amult25_Cmult61} {iopath_Amult25_Cmult62} {iopath_Amult25_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult26_Cmult26} {iopath_Amult26_Cmult27} {iopath_Amult26_Cmult28} {iopath_Amult26_Cmult29} {iopath_Amult26_Cmult30} {iopath_Amult26_Cmult31} {iopath_Amult26_Cmult32} {iopath_Amult26_Cmult33} {iopath_Amult26_Cmult34} {iopath_Amult26_Cmult35} {iopath_Amult26_Cmult36} {iopath_Amult26_Cmult37} {iopath_Amult26_Cmult38} {iopath_Amult26_Cmult39} {iopath_Amult26_Cmult40} {iopath_Amult26_Cmult41} {iopath_Amult26_Cmult42} {iopath_Amult26_Cmult43} {iopath_Amult26_Cmult44} {iopath_Amult26_Cmult45} {iopath_Amult26_Cmult46} {iopath_Amult26_Cmult47} {iopath_Amult26_Cmult48} {iopath_Amult26_Cmult49} {iopath_Amult26_Cmult50} {iopath_Amult26_Cmult51} {iopath_Amult26_Cmult52} {iopath_Amult26_Cmult53} {iopath_Amult26_Cmult54} {iopath_Amult26_Cmult55} {iopath_Amult26_Cmult56} {iopath_Amult26_Cmult57} {iopath_Amult26_Cmult58} {iopath_Amult26_Cmult59} {iopath_Amult26_Cmult60} {iopath_Amult26_Cmult61} {iopath_Amult26_Cmult62} {iopath_Amult26_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult27_Cmult27} {iopath_Amult27_Cmult28} {iopath_Amult27_Cmult29} {iopath_Amult27_Cmult30} {iopath_Amult27_Cmult31} {iopath_Amult27_Cmult32} {iopath_Amult27_Cmult33} {iopath_Amult27_Cmult34} {iopath_Amult27_Cmult35} {iopath_Amult27_Cmult36} {iopath_Amult27_Cmult37} {iopath_Amult27_Cmult38} {iopath_Amult27_Cmult39} {iopath_Amult27_Cmult40} {iopath_Amult27_Cmult41} {iopath_Amult27_Cmult42} {iopath_Amult27_Cmult43} {iopath_Amult27_Cmult44} {iopath_Amult27_Cmult45} {iopath_Amult27_Cmult46} {iopath_Amult27_Cmult47} {iopath_Amult27_Cmult48} {iopath_Amult27_Cmult49} {iopath_Amult27_Cmult50} {iopath_Amult27_Cmult51} {iopath_Amult27_Cmult52} {iopath_Amult27_Cmult53} {iopath_Amult27_Cmult54} {iopath_Amult27_Cmult55} {iopath_Amult27_Cmult56} {iopath_Amult27_Cmult57} {iopath_Amult27_Cmult58} {iopath_Amult27_Cmult59} {iopath_Amult27_Cmult60} {iopath_Amult27_Cmult61} {iopath_Amult27_Cmult62} {iopath_Amult27_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult28_Cmult28} {iopath_Amult28_Cmult29} {iopath_Amult28_Cmult30} {iopath_Amult28_Cmult31} {iopath_Amult28_Cmult32} {iopath_Amult28_Cmult33} {iopath_Amult28_Cmult34} {iopath_Amult28_Cmult35} {iopath_Amult28_Cmult36} {iopath_Amult28_Cmult37} {iopath_Amult28_Cmult38} {iopath_Amult28_Cmult39} {iopath_Amult28_Cmult40} {iopath_Amult28_Cmult41} {iopath_Amult28_Cmult42} {iopath_Amult28_Cmult43} {iopath_Amult28_Cmult44} {iopath_Amult28_Cmult45} {iopath_Amult28_Cmult46} {iopath_Amult28_Cmult47} {iopath_Amult28_Cmult48} {iopath_Amult28_Cmult49} {iopath_Amult28_Cmult50} {iopath_Amult28_Cmult51} {iopath_Amult28_Cmult52} {iopath_Amult28_Cmult53} {iopath_Amult28_Cmult54} {iopath_Amult28_Cmult55} {iopath_Amult28_Cmult56} {iopath_Amult28_Cmult57} {iopath_Amult28_Cmult58} {iopath_Amult28_Cmult59} {iopath_Amult28_Cmult60} {iopath_Amult28_Cmult61} {iopath_Amult28_Cmult62} {iopath_Amult28_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult29_Cmult29} {iopath_Amult29_Cmult30} {iopath_Amult29_Cmult31} {iopath_Amult29_Cmult32} {iopath_Amult29_Cmult33} {iopath_Amult29_Cmult34} {iopath_Amult29_Cmult35} {iopath_Amult29_Cmult36} {iopath_Amult29_Cmult37} {iopath_Amult29_Cmult38} {iopath_Amult29_Cmult39} {iopath_Amult29_Cmult40} {iopath_Amult29_Cmult41} {iopath_Amult29_Cmult42} {iopath_Amult29_Cmult43} {iopath_Amult29_Cmult44} {iopath_Amult29_Cmult45} {iopath_Amult29_Cmult46} {iopath_Amult29_Cmult47} {iopath_Amult29_Cmult48} {iopath_Amult29_Cmult49} {iopath_Amult29_Cmult50} {iopath_Amult29_Cmult51} {iopath_Amult29_Cmult52} {iopath_Amult29_Cmult53} {iopath_Amult29_Cmult54} {iopath_Amult29_Cmult55} {iopath_Amult29_Cmult56} {iopath_Amult29_Cmult57} {iopath_Amult29_Cmult58} {iopath_Amult29_Cmult59} {iopath_Amult29_Cmult60} {iopath_Amult29_Cmult61} {iopath_Amult29_Cmult62} {iopath_Amult29_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult30_Cmult30} {iopath_Amult30_Cmult31} {iopath_Amult30_Cmult32} {iopath_Amult30_Cmult33} {iopath_Amult30_Cmult34} {iopath_Amult30_Cmult35} {iopath_Amult30_Cmult36} {iopath_Amult30_Cmult37} {iopath_Amult30_Cmult38} {iopath_Amult30_Cmult39} {iopath_Amult30_Cmult40} {iopath_Amult30_Cmult41} {iopath_Amult30_Cmult42} {iopath_Amult30_Cmult43} {iopath_Amult30_Cmult44} {iopath_Amult30_Cmult45} {iopath_Amult30_Cmult46} {iopath_Amult30_Cmult47} {iopath_Amult30_Cmult48} {iopath_Amult30_Cmult49} {iopath_Amult30_Cmult50} {iopath_Amult30_Cmult51} {iopath_Amult30_Cmult52} {iopath_Amult30_Cmult53} {iopath_Amult30_Cmult54} {iopath_Amult30_Cmult55} {iopath_Amult30_Cmult56} {iopath_Amult30_Cmult57} {iopath_Amult30_Cmult58} {iopath_Amult30_Cmult59} {iopath_Amult30_Cmult60} {iopath_Amult30_Cmult61} {iopath_Amult30_Cmult62} {iopath_Amult30_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult31_Cmult31} {iopath_Amult31_Cmult32} {iopath_Amult31_Cmult33} {iopath_Amult31_Cmult34} {iopath_Amult31_Cmult35} {iopath_Amult31_Cmult36} {iopath_Amult31_Cmult37} {iopath_Amult31_Cmult38} {iopath_Amult31_Cmult39} {iopath_Amult31_Cmult40} {iopath_Amult31_Cmult41} {iopath_Amult31_Cmult42} {iopath_Amult31_Cmult43} {iopath_Amult31_Cmult44} {iopath_Amult31_Cmult45} {iopath_Amult31_Cmult46} {iopath_Amult31_Cmult47} {iopath_Amult31_Cmult48} {iopath_Amult31_Cmult49} {iopath_Amult31_Cmult50} {iopath_Amult31_Cmult51} {iopath_Amult31_Cmult52} {iopath_Amult31_Cmult53} {iopath_Amult31_Cmult54} {iopath_Amult31_Cmult55} {iopath_Amult31_Cmult56} {iopath_Amult31_Cmult57} {iopath_Amult31_Cmult58} {iopath_Amult31_Cmult59} {iopath_Amult31_Cmult60} {iopath_Amult31_Cmult61} {iopath_Amult31_Cmult62} {iopath_Amult31_Cmult63} "*)
	(* DELAY_MATRIX_Bmult="{iopath_Amult0_Cmult0} {iopath_Amult0_Cmult1} {iopath_Amult0_Cmult2} {iopath_Amult0_Cmult3} {iopath_Amult0_Cmult4} {iopath_Amult0_Cmult5} {iopath_Amult0_Cmult6} {iopath_Amult0_Cmult7} {iopath_Amult0_Cmult8} {iopath_Amult0_Cmult9} {iopath_Amult0_Cmult10} {iopath_Amult0_Cmult11} {iopath_Amult0_Cmult12} {iopath_Amult0_Cmult13} {iopath_Amult0_Cmult14} {iopath_Amult0_Cmult15} {iopath_Amult0_Cmult16} {iopath_Amult0_Cmult17} {iopath_Amult0_Cmult18} {iopath_Amult0_Cmult19} {iopath_Amult0_Cmult20} {iopath_Amult0_Cmult21} {iopath_Amult0_Cmult22} {iopath_Amult0_Cmult23} {iopath_Amult0_Cmult24} {iopath_Amult0_Cmult25} {iopath_Amult0_Cmult26} {iopath_Amult0_Cmult27} {iopath_Amult0_Cmult28} {iopath_Amult0_Cmult29} {iopath_Amult0_Cmult30} {iopath_Amult0_Cmult31} {iopath_Amult0_Cmult32} {iopath_Amult0_Cmult33} {iopath_Amult0_Cmult34} {iopath_Amult0_Cmult35} {iopath_Amult0_Cmult36} {iopath_Amult0_Cmult37} {iopath_Amult0_Cmult38} {iopath_Amult0_Cmult39} {iopath_Amult0_Cmult40} {iopath_Amult0_Cmult41} {iopath_Amult0_Cmult42} {iopath_Amult0_Cmult43} {iopath_Amult0_Cmult44} {iopath_Amult0_Cmult45} {iopath_Amult0_Cmult46} {iopath_Amult0_Cmult47} {iopath_Amult0_Cmult48} {iopath_Amult0_Cmult49} {iopath_Amult0_Cmult50} {iopath_Amult0_Cmult51} {iopath_Amult0_Cmult52} {iopath_Amult0_Cmult53} {iopath_Amult0_Cmult54} {iopath_Amult0_Cmult55} {iopath_Amult0_Cmult56} {iopath_Amult0_Cmult57} {iopath_Amult0_Cmult58} {iopath_Amult0_Cmult59} {iopath_Amult0_Cmult60} {iopath_Amult0_Cmult61} {iopath_Amult0_Cmult62} {iopath_Amult0_Cmult63} 0 {iopath_Amult1_Cmult1} {iopath_Amult1_Cmult2} {iopath_Amult1_Cmult3} {iopath_Amult1_Cmult4} {iopath_Amult1_Cmult5} {iopath_Amult1_Cmult6} {iopath_Amult1_Cmult7} {iopath_Amult1_Cmult8} {iopath_Amult1_Cmult9} {iopath_Amult1_Cmult10} {iopath_Amult1_Cmult11} {iopath_Amult1_Cmult12} {iopath_Amult1_Cmult13} {iopath_Amult1_Cmult14} {iopath_Amult1_Cmult15} {iopath_Amult1_Cmult16} {iopath_Amult1_Cmult17} {iopath_Amult1_Cmult18} {iopath_Amult1_Cmult19} {iopath_Amult1_Cmult20} {iopath_Amult1_Cmult21} {iopath_Amult1_Cmult22} {iopath_Amult1_Cmult23} {iopath_Amult1_Cmult24} {iopath_Amult1_Cmult25} {iopath_Amult1_Cmult26} {iopath_Amult1_Cmult27} {iopath_Amult1_Cmult28} {iopath_Amult1_Cmult29} {iopath_Amult1_Cmult30} {iopath_Amult1_Cmult31} {iopath_Amult1_Cmult32} {iopath_Amult1_Cmult33} {iopath_Amult1_Cmult34} {iopath_Amult1_Cmult35} {iopath_Amult1_Cmult36} {iopath_Amult1_Cmult37} {iopath_Amult1_Cmult38} {iopath_Amult1_Cmult39} {iopath_Amult1_Cmult40} {iopath_Amult1_Cmult41} {iopath_Amult1_Cmult42} {iopath_Amult1_Cmult43} {iopath_Amult1_Cmult44} {iopath_Amult1_Cmult45} {iopath_Amult1_Cmult46} {iopath_Amult1_Cmult47} {iopath_Amult1_Cmult48} {iopath_Amult1_Cmult49} {iopath_Amult1_Cmult50} {iopath_Amult1_Cmult51} {iopath_Amult1_Cmult52} {iopath_Amult1_Cmult53} {iopath_Amult1_Cmult54} {iopath_Amult1_Cmult55} {iopath_Amult1_Cmult56} {iopath_Amult1_Cmult57} {iopath_Amult1_Cmult58} {iopath_Amult1_Cmult59} {iopath_Amult1_Cmult60} {iopath_Amult1_Cmult61} {iopath_Amult1_Cmult62} {iopath_Amult1_Cmult63} 0 0 {iopath_Amult2_Cmult2} {iopath_Amult2_Cmult3} {iopath_Amult2_Cmult4} {iopath_Amult2_Cmult5} {iopath_Amult2_Cmult6} {iopath_Amult2_Cmult7} {iopath_Amult2_Cmult8} {iopath_Amult2_Cmult9} {iopath_Amult2_Cmult10} {iopath_Amult2_Cmult11} {iopath_Amult2_Cmult12} {iopath_Amult2_Cmult13} {iopath_Amult2_Cmult14} {iopath_Amult2_Cmult15} {iopath_Amult2_Cmult16} {iopath_Amult2_Cmult17} {iopath_Amult2_Cmult18} {iopath_Amult2_Cmult19} {iopath_Amult2_Cmult20} {iopath_Amult2_Cmult21} {iopath_Amult2_Cmult22} {iopath_Amult2_Cmult23} {iopath_Amult2_Cmult24} {iopath_Amult2_Cmult25} {iopath_Amult2_Cmult26} {iopath_Amult2_Cmult27} {iopath_Amult2_Cmult28} {iopath_Amult2_Cmult29} {iopath_Amult2_Cmult30} {iopath_Amult2_Cmult31} {iopath_Amult2_Cmult32} {iopath_Amult2_Cmult33} {iopath_Amult2_Cmult34} {iopath_Amult2_Cmult35} {iopath_Amult2_Cmult36} {iopath_Amult2_Cmult37} {iopath_Amult2_Cmult38} {iopath_Amult2_Cmult39} {iopath_Amult2_Cmult40} {iopath_Amult2_Cmult41} {iopath_Amult2_Cmult42} {iopath_Amult2_Cmult43} {iopath_Amult2_Cmult44} {iopath_Amult2_Cmult45} {iopath_Amult2_Cmult46} {iopath_Amult2_Cmult47} {iopath_Amult2_Cmult48} {iopath_Amult2_Cmult49} {iopath_Amult2_Cmult50} {iopath_Amult2_Cmult51} {iopath_Amult2_Cmult52} {iopath_Amult2_Cmult53} {iopath_Amult2_Cmult54} {iopath_Amult2_Cmult55} {iopath_Amult2_Cmult56} {iopath_Amult2_Cmult57} {iopath_Amult2_Cmult58} {iopath_Amult2_Cmult59} {iopath_Amult2_Cmult60} {iopath_Amult2_Cmult61} {iopath_Amult2_Cmult62} {iopath_Amult2_Cmult63} 0 0 0 {iopath_Amult3_Cmult3} {iopath_Amult3_Cmult4} {iopath_Amult3_Cmult5} {iopath_Amult3_Cmult6} {iopath_Amult3_Cmult7} {iopath_Amult3_Cmult8} {iopath_Amult3_Cmult9} {iopath_Amult3_Cmult10} {iopath_Amult3_Cmult11} {iopath_Amult3_Cmult12} {iopath_Amult3_Cmult13} {iopath_Amult3_Cmult14} {iopath_Amult3_Cmult15} {iopath_Amult3_Cmult16} {iopath_Amult3_Cmult17} {iopath_Amult3_Cmult18} {iopath_Amult3_Cmult19} {iopath_Amult3_Cmult20} {iopath_Amult3_Cmult21} {iopath_Amult3_Cmult22} {iopath_Amult3_Cmult23} {iopath_Amult3_Cmult24} {iopath_Amult3_Cmult25} {iopath_Amult3_Cmult26} {iopath_Amult3_Cmult27} {iopath_Amult3_Cmult28} {iopath_Amult3_Cmult29} {iopath_Amult3_Cmult30} {iopath_Amult3_Cmult31} {iopath_Amult3_Cmult32} {iopath_Amult3_Cmult33} {iopath_Amult3_Cmult34} {iopath_Amult3_Cmult35} {iopath_Amult3_Cmult36} {iopath_Amult3_Cmult37} {iopath_Amult3_Cmult38} {iopath_Amult3_Cmult39} {iopath_Amult3_Cmult40} {iopath_Amult3_Cmult41} {iopath_Amult3_Cmult42} {iopath_Amult3_Cmult43} {iopath_Amult3_Cmult44} {iopath_Amult3_Cmult45} {iopath_Amult3_Cmult46} {iopath_Amult3_Cmult47} {iopath_Amult3_Cmult48} {iopath_Amult3_Cmult49} {iopath_Amult3_Cmult50} {iopath_Amult3_Cmult51} {iopath_Amult3_Cmult52} {iopath_Amult3_Cmult53} {iopath_Amult3_Cmult54} {iopath_Amult3_Cmult55} {iopath_Amult3_Cmult56} {iopath_Amult3_Cmult57} {iopath_Amult3_Cmult58} {iopath_Amult3_Cmult59} {iopath_Amult3_Cmult60} {iopath_Amult3_Cmult61} {iopath_Amult3_Cmult62} {iopath_Amult3_Cmult63} 0 0 0 0 {iopath_Amult4_Cmult4} {iopath_Amult4_Cmult5} {iopath_Amult4_Cmult6} {iopath_Amult4_Cmult7} {iopath_Amult4_Cmult8} {iopath_Amult4_Cmult9} {iopath_Amult4_Cmult10} {iopath_Amult4_Cmult11} {iopath_Amult4_Cmult12} {iopath_Amult4_Cmult13} {iopath_Amult4_Cmult14} {iopath_Amult4_Cmult15} {iopath_Amult4_Cmult16} {iopath_Amult4_Cmult17} {iopath_Amult4_Cmult18} {iopath_Amult4_Cmult19} {iopath_Amult4_Cmult20} {iopath_Amult4_Cmult21} {iopath_Amult4_Cmult22} {iopath_Amult4_Cmult23} {iopath_Amult4_Cmult24} {iopath_Amult4_Cmult25} {iopath_Amult4_Cmult26} {iopath_Amult4_Cmult27} {iopath_Amult4_Cmult28} {iopath_Amult4_Cmult29} {iopath_Amult4_Cmult30} {iopath_Amult4_Cmult31} {iopath_Amult4_Cmult32} {iopath_Amult4_Cmult33} {iopath_Amult4_Cmult34} {iopath_Amult4_Cmult35} {iopath_Amult4_Cmult36} {iopath_Amult4_Cmult37} {iopath_Amult4_Cmult38} {iopath_Amult4_Cmult39} {iopath_Amult4_Cmult40} {iopath_Amult4_Cmult41} {iopath_Amult4_Cmult42} {iopath_Amult4_Cmult43} {iopath_Amult4_Cmult44} {iopath_Amult4_Cmult45} {iopath_Amult4_Cmult46} {iopath_Amult4_Cmult47} {iopath_Amult4_Cmult48} {iopath_Amult4_Cmult49} {iopath_Amult4_Cmult50} {iopath_Amult4_Cmult51} {iopath_Amult4_Cmult52} {iopath_Amult4_Cmult53} {iopath_Amult4_Cmult54} {iopath_Amult4_Cmult55} {iopath_Amult4_Cmult56} {iopath_Amult4_Cmult57} {iopath_Amult4_Cmult58} {iopath_Amult4_Cmult59} {iopath_Amult4_Cmult60} {iopath_Amult4_Cmult61} {iopath_Amult4_Cmult62} {iopath_Amult4_Cmult63} 0 0 0 0 0 {iopath_Amult5_Cmult5} {iopath_Amult5_Cmult6} {iopath_Amult5_Cmult7} {iopath_Amult5_Cmult8} {iopath_Amult5_Cmult9} {iopath_Amult5_Cmult10} {iopath_Amult5_Cmult11} {iopath_Amult5_Cmult12} {iopath_Amult5_Cmult13} {iopath_Amult5_Cmult14} {iopath_Amult5_Cmult15} {iopath_Amult5_Cmult16} {iopath_Amult5_Cmult17} {iopath_Amult5_Cmult18} {iopath_Amult5_Cmult19} {iopath_Amult5_Cmult20} {iopath_Amult5_Cmult21} {iopath_Amult5_Cmult22} {iopath_Amult5_Cmult23} {iopath_Amult5_Cmult24} {iopath_Amult5_Cmult25} {iopath_Amult5_Cmult26} {iopath_Amult5_Cmult27} {iopath_Amult5_Cmult28} {iopath_Amult5_Cmult29} {iopath_Amult5_Cmult30} {iopath_Amult5_Cmult31} {iopath_Amult5_Cmult32} {iopath_Amult5_Cmult33} {iopath_Amult5_Cmult34} {iopath_Amult5_Cmult35} {iopath_Amult5_Cmult36} {iopath_Amult5_Cmult37} {iopath_Amult5_Cmult38} {iopath_Amult5_Cmult39} {iopath_Amult5_Cmult40} {iopath_Amult5_Cmult41} {iopath_Amult5_Cmult42} {iopath_Amult5_Cmult43} {iopath_Amult5_Cmult44} {iopath_Amult5_Cmult45} {iopath_Amult5_Cmult46} {iopath_Amult5_Cmult47} {iopath_Amult5_Cmult48} {iopath_Amult5_Cmult49} {iopath_Amult5_Cmult50} {iopath_Amult5_Cmult51} {iopath_Amult5_Cmult52} {iopath_Amult5_Cmult53} {iopath_Amult5_Cmult54} {iopath_Amult5_Cmult55} {iopath_Amult5_Cmult56} {iopath_Amult5_Cmult57} {iopath_Amult5_Cmult58} {iopath_Amult5_Cmult59} {iopath_Amult5_Cmult60} {iopath_Amult5_Cmult61} {iopath_Amult5_Cmult62} {iopath_Amult5_Cmult63} 0 0 0 0 0 0 {iopath_Amult6_Cmult6} {iopath_Amult6_Cmult7} {iopath_Amult6_Cmult8} {iopath_Amult6_Cmult9} {iopath_Amult6_Cmult10} {iopath_Amult6_Cmult11} {iopath_Amult6_Cmult12} {iopath_Amult6_Cmult13} {iopath_Amult6_Cmult14} {iopath_Amult6_Cmult15} {iopath_Amult6_Cmult16} {iopath_Amult6_Cmult17} {iopath_Amult6_Cmult18} {iopath_Amult6_Cmult19} {iopath_Amult6_Cmult20} {iopath_Amult6_Cmult21} {iopath_Amult6_Cmult22} {iopath_Amult6_Cmult23} {iopath_Amult6_Cmult24} {iopath_Amult6_Cmult25} {iopath_Amult6_Cmult26} {iopath_Amult6_Cmult27} {iopath_Amult6_Cmult28} {iopath_Amult6_Cmult29} {iopath_Amult6_Cmult30} {iopath_Amult6_Cmult31} {iopath_Amult6_Cmult32} {iopath_Amult6_Cmult33} {iopath_Amult6_Cmult34} {iopath_Amult6_Cmult35} {iopath_Amult6_Cmult36} {iopath_Amult6_Cmult37} {iopath_Amult6_Cmult38} {iopath_Amult6_Cmult39} {iopath_Amult6_Cmult40} {iopath_Amult6_Cmult41} {iopath_Amult6_Cmult42} {iopath_Amult6_Cmult43} {iopath_Amult6_Cmult44} {iopath_Amult6_Cmult45} {iopath_Amult6_Cmult46} {iopath_Amult6_Cmult47} {iopath_Amult6_Cmult48} {iopath_Amult6_Cmult49} {iopath_Amult6_Cmult50} {iopath_Amult6_Cmult51} {iopath_Amult6_Cmult52} {iopath_Amult6_Cmult53} {iopath_Amult6_Cmult54} {iopath_Amult6_Cmult55} {iopath_Amult6_Cmult56} {iopath_Amult6_Cmult57} {iopath_Amult6_Cmult58} {iopath_Amult6_Cmult59} {iopath_Amult6_Cmult60} {iopath_Amult6_Cmult61} {iopath_Amult6_Cmult62} {iopath_Amult6_Cmult63} 0 0 0 0 0 0 0 {iopath_Amult7_Cmult7} {iopath_Amult7_Cmult8} {iopath_Amult7_Cmult9} {iopath_Amult7_Cmult10} {iopath_Amult7_Cmult11} {iopath_Amult7_Cmult12} {iopath_Amult7_Cmult13} {iopath_Amult7_Cmult14} {iopath_Amult7_Cmult15} {iopath_Amult7_Cmult16} {iopath_Amult7_Cmult17} {iopath_Amult7_Cmult18} {iopath_Amult7_Cmult19} {iopath_Amult7_Cmult20} {iopath_Amult7_Cmult21} {iopath_Amult7_Cmult22} {iopath_Amult7_Cmult23} {iopath_Amult7_Cmult24} {iopath_Amult7_Cmult25} {iopath_Amult7_Cmult26} {iopath_Amult7_Cmult27} {iopath_Amult7_Cmult28} {iopath_Amult7_Cmult29} {iopath_Amult7_Cmult30} {iopath_Amult7_Cmult31} {iopath_Amult7_Cmult32} {iopath_Amult7_Cmult33} {iopath_Amult7_Cmult34} {iopath_Amult7_Cmult35} {iopath_Amult7_Cmult36} {iopath_Amult7_Cmult37} {iopath_Amult7_Cmult38} {iopath_Amult7_Cmult39} {iopath_Amult7_Cmult40} {iopath_Amult7_Cmult41} {iopath_Amult7_Cmult42} {iopath_Amult7_Cmult43} {iopath_Amult7_Cmult44} {iopath_Amult7_Cmult45} {iopath_Amult7_Cmult46} {iopath_Amult7_Cmult47} {iopath_Amult7_Cmult48} {iopath_Amult7_Cmult49} {iopath_Amult7_Cmult50} {iopath_Amult7_Cmult51} {iopath_Amult7_Cmult52} {iopath_Amult7_Cmult53} {iopath_Amult7_Cmult54} {iopath_Amult7_Cmult55} {iopath_Amult7_Cmult56} {iopath_Amult7_Cmult57} {iopath_Amult7_Cmult58} {iopath_Amult7_Cmult59} {iopath_Amult7_Cmult60} {iopath_Amult7_Cmult61} {iopath_Amult7_Cmult62} {iopath_Amult7_Cmult63} 0 0 0 0 0 0 0 0 {iopath_Amult8_Cmult8} {iopath_Amult8_Cmult9} {iopath_Amult8_Cmult10} {iopath_Amult8_Cmult11} {iopath_Amult8_Cmult12} {iopath_Amult8_Cmult13} {iopath_Amult8_Cmult14} {iopath_Amult8_Cmult15} {iopath_Amult8_Cmult16} {iopath_Amult8_Cmult17} {iopath_Amult8_Cmult18} {iopath_Amult8_Cmult19} {iopath_Amult8_Cmult20} {iopath_Amult8_Cmult21} {iopath_Amult8_Cmult22} {iopath_Amult8_Cmult23} {iopath_Amult8_Cmult24} {iopath_Amult8_Cmult25} {iopath_Amult8_Cmult26} {iopath_Amult8_Cmult27} {iopath_Amult8_Cmult28} {iopath_Amult8_Cmult29} {iopath_Amult8_Cmult30} {iopath_Amult8_Cmult31} {iopath_Amult8_Cmult32} {iopath_Amult8_Cmult33} {iopath_Amult8_Cmult34} {iopath_Amult8_Cmult35} {iopath_Amult8_Cmult36} {iopath_Amult8_Cmult37} {iopath_Amult8_Cmult38} {iopath_Amult8_Cmult39} {iopath_Amult8_Cmult40} {iopath_Amult8_Cmult41} {iopath_Amult8_Cmult42} {iopath_Amult8_Cmult43} {iopath_Amult8_Cmult44} {iopath_Amult8_Cmult45} {iopath_Amult8_Cmult46} {iopath_Amult8_Cmult47} {iopath_Amult8_Cmult48} {iopath_Amult8_Cmult49} {iopath_Amult8_Cmult50} {iopath_Amult8_Cmult51} {iopath_Amult8_Cmult52} {iopath_Amult8_Cmult53} {iopath_Amult8_Cmult54} {iopath_Amult8_Cmult55} {iopath_Amult8_Cmult56} {iopath_Amult8_Cmult57} {iopath_Amult8_Cmult58} {iopath_Amult8_Cmult59} {iopath_Amult8_Cmult60} {iopath_Amult8_Cmult61} {iopath_Amult8_Cmult62} {iopath_Amult8_Cmult63} 0 0 0 0 0 0 0 0 0 {iopath_Amult9_Cmult9} {iopath_Amult9_Cmult10} {iopath_Amult9_Cmult11} {iopath_Amult9_Cmult12} {iopath_Amult9_Cmult13} {iopath_Amult9_Cmult14} {iopath_Amult9_Cmult15} {iopath_Amult9_Cmult16} {iopath_Amult9_Cmult17} {iopath_Amult9_Cmult18} {iopath_Amult9_Cmult19} {iopath_Amult9_Cmult20} {iopath_Amult9_Cmult21} {iopath_Amult9_Cmult22} {iopath_Amult9_Cmult23} {iopath_Amult9_Cmult24} {iopath_Amult9_Cmult25} {iopath_Amult9_Cmult26} {iopath_Amult9_Cmult27} {iopath_Amult9_Cmult28} {iopath_Amult9_Cmult29} {iopath_Amult9_Cmult30} {iopath_Amult9_Cmult31} {iopath_Amult9_Cmult32} {iopath_Amult9_Cmult33} {iopath_Amult9_Cmult34} {iopath_Amult9_Cmult35} {iopath_Amult9_Cmult36} {iopath_Amult9_Cmult37} {iopath_Amult9_Cmult38} {iopath_Amult9_Cmult39} {iopath_Amult9_Cmult40} {iopath_Amult9_Cmult41} {iopath_Amult9_Cmult42} {iopath_Amult9_Cmult43} {iopath_Amult9_Cmult44} {iopath_Amult9_Cmult45} {iopath_Amult9_Cmult46} {iopath_Amult9_Cmult47} {iopath_Amult9_Cmult48} {iopath_Amult9_Cmult49} {iopath_Amult9_Cmult50} {iopath_Amult9_Cmult51} {iopath_Amult9_Cmult52} {iopath_Amult9_Cmult53} {iopath_Amult9_Cmult54} {iopath_Amult9_Cmult55} {iopath_Amult9_Cmult56} {iopath_Amult9_Cmult57} {iopath_Amult9_Cmult58} {iopath_Amult9_Cmult59} {iopath_Amult9_Cmult60} {iopath_Amult9_Cmult61} {iopath_Amult9_Cmult62} {iopath_Amult9_Cmult63} 0 0 0 0 0 0 0 0 0 0 {iopath_Amult10_Cmult10} {iopath_Amult10_Cmult11} {iopath_Amult10_Cmult12} {iopath_Amult10_Cmult13} {iopath_Amult10_Cmult14} {iopath_Amult10_Cmult15} {iopath_Amult10_Cmult16} {iopath_Amult10_Cmult17} {iopath_Amult10_Cmult18} {iopath_Amult10_Cmult19} {iopath_Amult10_Cmult20} {iopath_Amult10_Cmult21} {iopath_Amult10_Cmult22} {iopath_Amult10_Cmult23} {iopath_Amult10_Cmult24} {iopath_Amult10_Cmult25} {iopath_Amult10_Cmult26} {iopath_Amult10_Cmult27} {iopath_Amult10_Cmult28} {iopath_Amult10_Cmult29} {iopath_Amult10_Cmult30} {iopath_Amult10_Cmult31} {iopath_Amult10_Cmult32} {iopath_Amult10_Cmult33} {iopath_Amult10_Cmult34} {iopath_Amult10_Cmult35} {iopath_Amult10_Cmult36} {iopath_Amult10_Cmult37} {iopath_Amult10_Cmult38} {iopath_Amult10_Cmult39} {iopath_Amult10_Cmult40} {iopath_Amult10_Cmult41} {iopath_Amult10_Cmult42} {iopath_Amult10_Cmult43} {iopath_Amult10_Cmult44} {iopath_Amult10_Cmult45} {iopath_Amult10_Cmult46} {iopath_Amult10_Cmult47} {iopath_Amult10_Cmult48} {iopath_Amult10_Cmult49} {iopath_Amult10_Cmult50} {iopath_Amult10_Cmult51} {iopath_Amult10_Cmult52} {iopath_Amult10_Cmult53} {iopath_Amult10_Cmult54} {iopath_Amult10_Cmult55} {iopath_Amult10_Cmult56} {iopath_Amult10_Cmult57} {iopath_Amult10_Cmult58} {iopath_Amult10_Cmult59} {iopath_Amult10_Cmult60} {iopath_Amult10_Cmult61} {iopath_Amult10_Cmult62} {iopath_Amult10_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult11_Cmult11} {iopath_Amult11_Cmult12} {iopath_Amult11_Cmult13} {iopath_Amult11_Cmult14} {iopath_Amult11_Cmult15} {iopath_Amult11_Cmult16} {iopath_Amult11_Cmult17} {iopath_Amult11_Cmult18} {iopath_Amult11_Cmult19} {iopath_Amult11_Cmult20} {iopath_Amult11_Cmult21} {iopath_Amult11_Cmult22} {iopath_Amult11_Cmult23} {iopath_Amult11_Cmult24} {iopath_Amult11_Cmult25} {iopath_Amult11_Cmult26} {iopath_Amult11_Cmult27} {iopath_Amult11_Cmult28} {iopath_Amult11_Cmult29} {iopath_Amult11_Cmult30} {iopath_Amult11_Cmult31} {iopath_Amult11_Cmult32} {iopath_Amult11_Cmult33} {iopath_Amult11_Cmult34} {iopath_Amult11_Cmult35} {iopath_Amult11_Cmult36} {iopath_Amult11_Cmult37} {iopath_Amult11_Cmult38} {iopath_Amult11_Cmult39} {iopath_Amult11_Cmult40} {iopath_Amult11_Cmult41} {iopath_Amult11_Cmult42} {iopath_Amult11_Cmult43} {iopath_Amult11_Cmult44} {iopath_Amult11_Cmult45} {iopath_Amult11_Cmult46} {iopath_Amult11_Cmult47} {iopath_Amult11_Cmult48} {iopath_Amult11_Cmult49} {iopath_Amult11_Cmult50} {iopath_Amult11_Cmult51} {iopath_Amult11_Cmult52} {iopath_Amult11_Cmult53} {iopath_Amult11_Cmult54} {iopath_Amult11_Cmult55} {iopath_Amult11_Cmult56} {iopath_Amult11_Cmult57} {iopath_Amult11_Cmult58} {iopath_Amult11_Cmult59} {iopath_Amult11_Cmult60} {iopath_Amult11_Cmult61} {iopath_Amult11_Cmult62} {iopath_Amult11_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult12_Cmult12} {iopath_Amult12_Cmult13} {iopath_Amult12_Cmult14} {iopath_Amult12_Cmult15} {iopath_Amult12_Cmult16} {iopath_Amult12_Cmult17} {iopath_Amult12_Cmult18} {iopath_Amult12_Cmult19} {iopath_Amult12_Cmult20} {iopath_Amult12_Cmult21} {iopath_Amult12_Cmult22} {iopath_Amult12_Cmult23} {iopath_Amult12_Cmult24} {iopath_Amult12_Cmult25} {iopath_Amult12_Cmult26} {iopath_Amult12_Cmult27} {iopath_Amult12_Cmult28} {iopath_Amult12_Cmult29} {iopath_Amult12_Cmult30} {iopath_Amult12_Cmult31} {iopath_Amult12_Cmult32} {iopath_Amult12_Cmult33} {iopath_Amult12_Cmult34} {iopath_Amult12_Cmult35} {iopath_Amult12_Cmult36} {iopath_Amult12_Cmult37} {iopath_Amult12_Cmult38} {iopath_Amult12_Cmult39} {iopath_Amult12_Cmult40} {iopath_Amult12_Cmult41} {iopath_Amult12_Cmult42} {iopath_Amult12_Cmult43} {iopath_Amult12_Cmult44} {iopath_Amult12_Cmult45} {iopath_Amult12_Cmult46} {iopath_Amult12_Cmult47} {iopath_Amult12_Cmult48} {iopath_Amult12_Cmult49} {iopath_Amult12_Cmult50} {iopath_Amult12_Cmult51} {iopath_Amult12_Cmult52} {iopath_Amult12_Cmult53} {iopath_Amult12_Cmult54} {iopath_Amult12_Cmult55} {iopath_Amult12_Cmult56} {iopath_Amult12_Cmult57} {iopath_Amult12_Cmult58} {iopath_Amult12_Cmult59} {iopath_Amult12_Cmult60} {iopath_Amult12_Cmult61} {iopath_Amult12_Cmult62} {iopath_Amult12_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult13_Cmult13} {iopath_Amult13_Cmult14} {iopath_Amult13_Cmult15} {iopath_Amult13_Cmult16} {iopath_Amult13_Cmult17} {iopath_Amult13_Cmult18} {iopath_Amult13_Cmult19} {iopath_Amult13_Cmult20} {iopath_Amult13_Cmult21} {iopath_Amult13_Cmult22} {iopath_Amult13_Cmult23} {iopath_Amult13_Cmult24} {iopath_Amult13_Cmult25} {iopath_Amult13_Cmult26} {iopath_Amult13_Cmult27} {iopath_Amult13_Cmult28} {iopath_Amult13_Cmult29} {iopath_Amult13_Cmult30} {iopath_Amult13_Cmult31} {iopath_Amult13_Cmult32} {iopath_Amult13_Cmult33} {iopath_Amult13_Cmult34} {iopath_Amult13_Cmult35} {iopath_Amult13_Cmult36} {iopath_Amult13_Cmult37} {iopath_Amult13_Cmult38} {iopath_Amult13_Cmult39} {iopath_Amult13_Cmult40} {iopath_Amult13_Cmult41} {iopath_Amult13_Cmult42} {iopath_Amult13_Cmult43} {iopath_Amult13_Cmult44} {iopath_Amult13_Cmult45} {iopath_Amult13_Cmult46} {iopath_Amult13_Cmult47} {iopath_Amult13_Cmult48} {iopath_Amult13_Cmult49} {iopath_Amult13_Cmult50} {iopath_Amult13_Cmult51} {iopath_Amult13_Cmult52} {iopath_Amult13_Cmult53} {iopath_Amult13_Cmult54} {iopath_Amult13_Cmult55} {iopath_Amult13_Cmult56} {iopath_Amult13_Cmult57} {iopath_Amult13_Cmult58} {iopath_Amult13_Cmult59} {iopath_Amult13_Cmult60} {iopath_Amult13_Cmult61} {iopath_Amult13_Cmult62} {iopath_Amult13_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult14_Cmult14} {iopath_Amult14_Cmult15} {iopath_Amult14_Cmult16} {iopath_Amult14_Cmult17} {iopath_Amult14_Cmult18} {iopath_Amult14_Cmult19} {iopath_Amult14_Cmult20} {iopath_Amult14_Cmult21} {iopath_Amult14_Cmult22} {iopath_Amult14_Cmult23} {iopath_Amult14_Cmult24} {iopath_Amult14_Cmult25} {iopath_Amult14_Cmult26} {iopath_Amult14_Cmult27} {iopath_Amult14_Cmult28} {iopath_Amult14_Cmult29} {iopath_Amult14_Cmult30} {iopath_Amult14_Cmult31} {iopath_Amult14_Cmult32} {iopath_Amult14_Cmult33} {iopath_Amult14_Cmult34} {iopath_Amult14_Cmult35} {iopath_Amult14_Cmult36} {iopath_Amult14_Cmult37} {iopath_Amult14_Cmult38} {iopath_Amult14_Cmult39} {iopath_Amult14_Cmult40} {iopath_Amult14_Cmult41} {iopath_Amult14_Cmult42} {iopath_Amult14_Cmult43} {iopath_Amult14_Cmult44} {iopath_Amult14_Cmult45} {iopath_Amult14_Cmult46} {iopath_Amult14_Cmult47} {iopath_Amult14_Cmult48} {iopath_Amult14_Cmult49} {iopath_Amult14_Cmult50} {iopath_Amult14_Cmult51} {iopath_Amult14_Cmult52} {iopath_Amult14_Cmult53} {iopath_Amult14_Cmult54} {iopath_Amult14_Cmult55} {iopath_Amult14_Cmult56} {iopath_Amult14_Cmult57} {iopath_Amult14_Cmult58} {iopath_Amult14_Cmult59} {iopath_Amult14_Cmult60} {iopath_Amult14_Cmult61} {iopath_Amult14_Cmult62} {iopath_Amult14_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult15_Cmult15} {iopath_Amult15_Cmult16} {iopath_Amult15_Cmult17} {iopath_Amult15_Cmult18} {iopath_Amult15_Cmult19} {iopath_Amult15_Cmult20} {iopath_Amult15_Cmult21} {iopath_Amult15_Cmult22} {iopath_Amult15_Cmult23} {iopath_Amult15_Cmult24} {iopath_Amult15_Cmult25} {iopath_Amult15_Cmult26} {iopath_Amult15_Cmult27} {iopath_Amult15_Cmult28} {iopath_Amult15_Cmult29} {iopath_Amult15_Cmult30} {iopath_Amult15_Cmult31} {iopath_Amult15_Cmult32} {iopath_Amult15_Cmult33} {iopath_Amult15_Cmult34} {iopath_Amult15_Cmult35} {iopath_Amult15_Cmult36} {iopath_Amult15_Cmult37} {iopath_Amult15_Cmult38} {iopath_Amult15_Cmult39} {iopath_Amult15_Cmult40} {iopath_Amult15_Cmult41} {iopath_Amult15_Cmult42} {iopath_Amult15_Cmult43} {iopath_Amult15_Cmult44} {iopath_Amult15_Cmult45} {iopath_Amult15_Cmult46} {iopath_Amult15_Cmult47} {iopath_Amult15_Cmult48} {iopath_Amult15_Cmult49} {iopath_Amult15_Cmult50} {iopath_Amult15_Cmult51} {iopath_Amult15_Cmult52} {iopath_Amult15_Cmult53} {iopath_Amult15_Cmult54} {iopath_Amult15_Cmult55} {iopath_Amult15_Cmult56} {iopath_Amult15_Cmult57} {iopath_Amult15_Cmult58} {iopath_Amult15_Cmult59} {iopath_Amult15_Cmult60} {iopath_Amult15_Cmult61} {iopath_Amult15_Cmult62} {iopath_Amult15_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult16_Cmult16} {iopath_Amult16_Cmult17} {iopath_Amult16_Cmult18} {iopath_Amult16_Cmult19} {iopath_Amult16_Cmult20} {iopath_Amult16_Cmult21} {iopath_Amult16_Cmult22} {iopath_Amult16_Cmult23} {iopath_Amult16_Cmult24} {iopath_Amult16_Cmult25} {iopath_Amult16_Cmult26} {iopath_Amult16_Cmult27} {iopath_Amult16_Cmult28} {iopath_Amult16_Cmult29} {iopath_Amult16_Cmult30} {iopath_Amult16_Cmult31} {iopath_Amult16_Cmult32} {iopath_Amult16_Cmult33} {iopath_Amult16_Cmult34} {iopath_Amult16_Cmult35} {iopath_Amult16_Cmult36} {iopath_Amult16_Cmult37} {iopath_Amult16_Cmult38} {iopath_Amult16_Cmult39} {iopath_Amult16_Cmult40} {iopath_Amult16_Cmult41} {iopath_Amult16_Cmult42} {iopath_Amult16_Cmult43} {iopath_Amult16_Cmult44} {iopath_Amult16_Cmult45} {iopath_Amult16_Cmult46} {iopath_Amult16_Cmult47} {iopath_Amult16_Cmult48} {iopath_Amult16_Cmult49} {iopath_Amult16_Cmult50} {iopath_Amult16_Cmult51} {iopath_Amult16_Cmult52} {iopath_Amult16_Cmult53} {iopath_Amult16_Cmult54} {iopath_Amult16_Cmult55} {iopath_Amult16_Cmult56} {iopath_Amult16_Cmult57} {iopath_Amult16_Cmult58} {iopath_Amult16_Cmult59} {iopath_Amult16_Cmult60} {iopath_Amult16_Cmult61} {iopath_Amult16_Cmult62} {iopath_Amult16_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult17_Cmult17} {iopath_Amult17_Cmult18} {iopath_Amult17_Cmult19} {iopath_Amult17_Cmult20} {iopath_Amult17_Cmult21} {iopath_Amult17_Cmult22} {iopath_Amult17_Cmult23} {iopath_Amult17_Cmult24} {iopath_Amult17_Cmult25} {iopath_Amult17_Cmult26} {iopath_Amult17_Cmult27} {iopath_Amult17_Cmult28} {iopath_Amult17_Cmult29} {iopath_Amult17_Cmult30} {iopath_Amult17_Cmult31} {iopath_Amult17_Cmult32} {iopath_Amult17_Cmult33} {iopath_Amult17_Cmult34} {iopath_Amult17_Cmult35} {iopath_Amult17_Cmult36} {iopath_Amult17_Cmult37} {iopath_Amult17_Cmult38} {iopath_Amult17_Cmult39} {iopath_Amult17_Cmult40} {iopath_Amult17_Cmult41} {iopath_Amult17_Cmult42} {iopath_Amult17_Cmult43} {iopath_Amult17_Cmult44} {iopath_Amult17_Cmult45} {iopath_Amult17_Cmult46} {iopath_Amult17_Cmult47} {iopath_Amult17_Cmult48} {iopath_Amult17_Cmult49} {iopath_Amult17_Cmult50} {iopath_Amult17_Cmult51} {iopath_Amult17_Cmult52} {iopath_Amult17_Cmult53} {iopath_Amult17_Cmult54} {iopath_Amult17_Cmult55} {iopath_Amult17_Cmult56} {iopath_Amult17_Cmult57} {iopath_Amult17_Cmult58} {iopath_Amult17_Cmult59} {iopath_Amult17_Cmult60} {iopath_Amult17_Cmult61} {iopath_Amult17_Cmult62} {iopath_Amult17_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult18_Cmult18} {iopath_Amult18_Cmult19} {iopath_Amult18_Cmult20} {iopath_Amult18_Cmult21} {iopath_Amult18_Cmult22} {iopath_Amult18_Cmult23} {iopath_Amult18_Cmult24} {iopath_Amult18_Cmult25} {iopath_Amult18_Cmult26} {iopath_Amult18_Cmult27} {iopath_Amult18_Cmult28} {iopath_Amult18_Cmult29} {iopath_Amult18_Cmult30} {iopath_Amult18_Cmult31} {iopath_Amult18_Cmult32} {iopath_Amult18_Cmult33} {iopath_Amult18_Cmult34} {iopath_Amult18_Cmult35} {iopath_Amult18_Cmult36} {iopath_Amult18_Cmult37} {iopath_Amult18_Cmult38} {iopath_Amult18_Cmult39} {iopath_Amult18_Cmult40} {iopath_Amult18_Cmult41} {iopath_Amult18_Cmult42} {iopath_Amult18_Cmult43} {iopath_Amult18_Cmult44} {iopath_Amult18_Cmult45} {iopath_Amult18_Cmult46} {iopath_Amult18_Cmult47} {iopath_Amult18_Cmult48} {iopath_Amult18_Cmult49} {iopath_Amult18_Cmult50} {iopath_Amult18_Cmult51} {iopath_Amult18_Cmult52} {iopath_Amult18_Cmult53} {iopath_Amult18_Cmult54} {iopath_Amult18_Cmult55} {iopath_Amult18_Cmult56} {iopath_Amult18_Cmult57} {iopath_Amult18_Cmult58} {iopath_Amult18_Cmult59} {iopath_Amult18_Cmult60} {iopath_Amult18_Cmult61} {iopath_Amult18_Cmult62} {iopath_Amult18_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult19_Cmult19} {iopath_Amult19_Cmult20} {iopath_Amult19_Cmult21} {iopath_Amult19_Cmult22} {iopath_Amult19_Cmult23} {iopath_Amult19_Cmult24} {iopath_Amult19_Cmult25} {iopath_Amult19_Cmult26} {iopath_Amult19_Cmult27} {iopath_Amult19_Cmult28} {iopath_Amult19_Cmult29} {iopath_Amult19_Cmult30} {iopath_Amult19_Cmult31} {iopath_Amult19_Cmult32} {iopath_Amult19_Cmult33} {iopath_Amult19_Cmult34} {iopath_Amult19_Cmult35} {iopath_Amult19_Cmult36} {iopath_Amult19_Cmult37} {iopath_Amult19_Cmult38} {iopath_Amult19_Cmult39} {iopath_Amult19_Cmult40} {iopath_Amult19_Cmult41} {iopath_Amult19_Cmult42} {iopath_Amult19_Cmult43} {iopath_Amult19_Cmult44} {iopath_Amult19_Cmult45} {iopath_Amult19_Cmult46} {iopath_Amult19_Cmult47} {iopath_Amult19_Cmult48} {iopath_Amult19_Cmult49} {iopath_Amult19_Cmult50} {iopath_Amult19_Cmult51} {iopath_Amult19_Cmult52} {iopath_Amult19_Cmult53} {iopath_Amult19_Cmult54} {iopath_Amult19_Cmult55} {iopath_Amult19_Cmult56} {iopath_Amult19_Cmult57} {iopath_Amult19_Cmult58} {iopath_Amult19_Cmult59} {iopath_Amult19_Cmult60} {iopath_Amult19_Cmult61} {iopath_Amult19_Cmult62} {iopath_Amult19_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult20_Cmult20} {iopath_Amult20_Cmult21} {iopath_Amult20_Cmult22} {iopath_Amult20_Cmult23} {iopath_Amult20_Cmult24} {iopath_Amult20_Cmult25} {iopath_Amult20_Cmult26} {iopath_Amult20_Cmult27} {iopath_Amult20_Cmult28} {iopath_Amult20_Cmult29} {iopath_Amult20_Cmult30} {iopath_Amult20_Cmult31} {iopath_Amult20_Cmult32} {iopath_Amult20_Cmult33} {iopath_Amult20_Cmult34} {iopath_Amult20_Cmult35} {iopath_Amult20_Cmult36} {iopath_Amult20_Cmult37} {iopath_Amult20_Cmult38} {iopath_Amult20_Cmult39} {iopath_Amult20_Cmult40} {iopath_Amult20_Cmult41} {iopath_Amult20_Cmult42} {iopath_Amult20_Cmult43} {iopath_Amult20_Cmult44} {iopath_Amult20_Cmult45} {iopath_Amult20_Cmult46} {iopath_Amult20_Cmult47} {iopath_Amult20_Cmult48} {iopath_Amult20_Cmult49} {iopath_Amult20_Cmult50} {iopath_Amult20_Cmult51} {iopath_Amult20_Cmult52} {iopath_Amult20_Cmult53} {iopath_Amult20_Cmult54} {iopath_Amult20_Cmult55} {iopath_Amult20_Cmult56} {iopath_Amult20_Cmult57} {iopath_Amult20_Cmult58} {iopath_Amult20_Cmult59} {iopath_Amult20_Cmult60} {iopath_Amult20_Cmult61} {iopath_Amult20_Cmult62} {iopath_Amult20_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult21_Cmult21} {iopath_Amult21_Cmult22} {iopath_Amult21_Cmult23} {iopath_Amult21_Cmult24} {iopath_Amult21_Cmult25} {iopath_Amult21_Cmult26} {iopath_Amult21_Cmult27} {iopath_Amult21_Cmult28} {iopath_Amult21_Cmult29} {iopath_Amult21_Cmult30} {iopath_Amult21_Cmult31} {iopath_Amult21_Cmult32} {iopath_Amult21_Cmult33} {iopath_Amult21_Cmult34} {iopath_Amult21_Cmult35} {iopath_Amult21_Cmult36} {iopath_Amult21_Cmult37} {iopath_Amult21_Cmult38} {iopath_Amult21_Cmult39} {iopath_Amult21_Cmult40} {iopath_Amult21_Cmult41} {iopath_Amult21_Cmult42} {iopath_Amult21_Cmult43} {iopath_Amult21_Cmult44} {iopath_Amult21_Cmult45} {iopath_Amult21_Cmult46} {iopath_Amult21_Cmult47} {iopath_Amult21_Cmult48} {iopath_Amult21_Cmult49} {iopath_Amult21_Cmult50} {iopath_Amult21_Cmult51} {iopath_Amult21_Cmult52} {iopath_Amult21_Cmult53} {iopath_Amult21_Cmult54} {iopath_Amult21_Cmult55} {iopath_Amult21_Cmult56} {iopath_Amult21_Cmult57} {iopath_Amult21_Cmult58} {iopath_Amult21_Cmult59} {iopath_Amult21_Cmult60} {iopath_Amult21_Cmult61} {iopath_Amult21_Cmult62} {iopath_Amult21_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult22_Cmult22} {iopath_Amult22_Cmult23} {iopath_Amult22_Cmult24} {iopath_Amult22_Cmult25} {iopath_Amult22_Cmult26} {iopath_Amult22_Cmult27} {iopath_Amult22_Cmult28} {iopath_Amult22_Cmult29} {iopath_Amult22_Cmult30} {iopath_Amult22_Cmult31} {iopath_Amult22_Cmult32} {iopath_Amult22_Cmult33} {iopath_Amult22_Cmult34} {iopath_Amult22_Cmult35} {iopath_Amult22_Cmult36} {iopath_Amult22_Cmult37} {iopath_Amult22_Cmult38} {iopath_Amult22_Cmult39} {iopath_Amult22_Cmult40} {iopath_Amult22_Cmult41} {iopath_Amult22_Cmult42} {iopath_Amult22_Cmult43} {iopath_Amult22_Cmult44} {iopath_Amult22_Cmult45} {iopath_Amult22_Cmult46} {iopath_Amult22_Cmult47} {iopath_Amult22_Cmult48} {iopath_Amult22_Cmult49} {iopath_Amult22_Cmult50} {iopath_Amult22_Cmult51} {iopath_Amult22_Cmult52} {iopath_Amult22_Cmult53} {iopath_Amult22_Cmult54} {iopath_Amult22_Cmult55} {iopath_Amult22_Cmult56} {iopath_Amult22_Cmult57} {iopath_Amult22_Cmult58} {iopath_Amult22_Cmult59} {iopath_Amult22_Cmult60} {iopath_Amult22_Cmult61} {iopath_Amult22_Cmult62} {iopath_Amult22_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult23_Cmult23} {iopath_Amult23_Cmult24} {iopath_Amult23_Cmult25} {iopath_Amult23_Cmult26} {iopath_Amult23_Cmult27} {iopath_Amult23_Cmult28} {iopath_Amult23_Cmult29} {iopath_Amult23_Cmult30} {iopath_Amult23_Cmult31} {iopath_Amult23_Cmult32} {iopath_Amult23_Cmult33} {iopath_Amult23_Cmult34} {iopath_Amult23_Cmult35} {iopath_Amult23_Cmult36} {iopath_Amult23_Cmult37} {iopath_Amult23_Cmult38} {iopath_Amult23_Cmult39} {iopath_Amult23_Cmult40} {iopath_Amult23_Cmult41} {iopath_Amult23_Cmult42} {iopath_Amult23_Cmult43} {iopath_Amult23_Cmult44} {iopath_Amult23_Cmult45} {iopath_Amult23_Cmult46} {iopath_Amult23_Cmult47} {iopath_Amult23_Cmult48} {iopath_Amult23_Cmult49} {iopath_Amult23_Cmult50} {iopath_Amult23_Cmult51} {iopath_Amult23_Cmult52} {iopath_Amult23_Cmult53} {iopath_Amult23_Cmult54} {iopath_Amult23_Cmult55} {iopath_Amult23_Cmult56} {iopath_Amult23_Cmult57} {iopath_Amult23_Cmult58} {iopath_Amult23_Cmult59} {iopath_Amult23_Cmult60} {iopath_Amult23_Cmult61} {iopath_Amult23_Cmult62} {iopath_Amult23_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult24_Cmult24} {iopath_Amult24_Cmult25} {iopath_Amult24_Cmult26} {iopath_Amult24_Cmult27} {iopath_Amult24_Cmult28} {iopath_Amult24_Cmult29} {iopath_Amult24_Cmult30} {iopath_Amult24_Cmult31} {iopath_Amult24_Cmult32} {iopath_Amult24_Cmult33} {iopath_Amult24_Cmult34} {iopath_Amult24_Cmult35} {iopath_Amult24_Cmult36} {iopath_Amult24_Cmult37} {iopath_Amult24_Cmult38} {iopath_Amult24_Cmult39} {iopath_Amult24_Cmult40} {iopath_Amult24_Cmult41} {iopath_Amult24_Cmult42} {iopath_Amult24_Cmult43} {iopath_Amult24_Cmult44} {iopath_Amult24_Cmult45} {iopath_Amult24_Cmult46} {iopath_Amult24_Cmult47} {iopath_Amult24_Cmult48} {iopath_Amult24_Cmult49} {iopath_Amult24_Cmult50} {iopath_Amult24_Cmult51} {iopath_Amult24_Cmult52} {iopath_Amult24_Cmult53} {iopath_Amult24_Cmult54} {iopath_Amult24_Cmult55} {iopath_Amult24_Cmult56} {iopath_Amult24_Cmult57} {iopath_Amult24_Cmult58} {iopath_Amult24_Cmult59} {iopath_Amult24_Cmult60} {iopath_Amult24_Cmult61} {iopath_Amult24_Cmult62} {iopath_Amult24_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult25_Cmult25} {iopath_Amult25_Cmult26} {iopath_Amult25_Cmult27} {iopath_Amult25_Cmult28} {iopath_Amult25_Cmult29} {iopath_Amult25_Cmult30} {iopath_Amult25_Cmult31} {iopath_Amult25_Cmult32} {iopath_Amult25_Cmult33} {iopath_Amult25_Cmult34} {iopath_Amult25_Cmult35} {iopath_Amult25_Cmult36} {iopath_Amult25_Cmult37} {iopath_Amult25_Cmult38} {iopath_Amult25_Cmult39} {iopath_Amult25_Cmult40} {iopath_Amult25_Cmult41} {iopath_Amult25_Cmult42} {iopath_Amult25_Cmult43} {iopath_Amult25_Cmult44} {iopath_Amult25_Cmult45} {iopath_Amult25_Cmult46} {iopath_Amult25_Cmult47} {iopath_Amult25_Cmult48} {iopath_Amult25_Cmult49} {iopath_Amult25_Cmult50} {iopath_Amult25_Cmult51} {iopath_Amult25_Cmult52} {iopath_Amult25_Cmult53} {iopath_Amult25_Cmult54} {iopath_Amult25_Cmult55} {iopath_Amult25_Cmult56} {iopath_Amult25_Cmult57} {iopath_Amult25_Cmult58} {iopath_Amult25_Cmult59} {iopath_Amult25_Cmult60} {iopath_Amult25_Cmult61} {iopath_Amult25_Cmult62} {iopath_Amult25_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult26_Cmult26} {iopath_Amult26_Cmult27} {iopath_Amult26_Cmult28} {iopath_Amult26_Cmult29} {iopath_Amult26_Cmult30} {iopath_Amult26_Cmult31} {iopath_Amult26_Cmult32} {iopath_Amult26_Cmult33} {iopath_Amult26_Cmult34} {iopath_Amult26_Cmult35} {iopath_Amult26_Cmult36} {iopath_Amult26_Cmult37} {iopath_Amult26_Cmult38} {iopath_Amult26_Cmult39} {iopath_Amult26_Cmult40} {iopath_Amult26_Cmult41} {iopath_Amult26_Cmult42} {iopath_Amult26_Cmult43} {iopath_Amult26_Cmult44} {iopath_Amult26_Cmult45} {iopath_Amult26_Cmult46} {iopath_Amult26_Cmult47} {iopath_Amult26_Cmult48} {iopath_Amult26_Cmult49} {iopath_Amult26_Cmult50} {iopath_Amult26_Cmult51} {iopath_Amult26_Cmult52} {iopath_Amult26_Cmult53} {iopath_Amult26_Cmult54} {iopath_Amult26_Cmult55} {iopath_Amult26_Cmult56} {iopath_Amult26_Cmult57} {iopath_Amult26_Cmult58} {iopath_Amult26_Cmult59} {iopath_Amult26_Cmult60} {iopath_Amult26_Cmult61} {iopath_Amult26_Cmult62} {iopath_Amult26_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult27_Cmult27} {iopath_Amult27_Cmult28} {iopath_Amult27_Cmult29} {iopath_Amult27_Cmult30} {iopath_Amult27_Cmult31} {iopath_Amult27_Cmult32} {iopath_Amult27_Cmult33} {iopath_Amult27_Cmult34} {iopath_Amult27_Cmult35} {iopath_Amult27_Cmult36} {iopath_Amult27_Cmult37} {iopath_Amult27_Cmult38} {iopath_Amult27_Cmult39} {iopath_Amult27_Cmult40} {iopath_Amult27_Cmult41} {iopath_Amult27_Cmult42} {iopath_Amult27_Cmult43} {iopath_Amult27_Cmult44} {iopath_Amult27_Cmult45} {iopath_Amult27_Cmult46} {iopath_Amult27_Cmult47} {iopath_Amult27_Cmult48} {iopath_Amult27_Cmult49} {iopath_Amult27_Cmult50} {iopath_Amult27_Cmult51} {iopath_Amult27_Cmult52} {iopath_Amult27_Cmult53} {iopath_Amult27_Cmult54} {iopath_Amult27_Cmult55} {iopath_Amult27_Cmult56} {iopath_Amult27_Cmult57} {iopath_Amult27_Cmult58} {iopath_Amult27_Cmult59} {iopath_Amult27_Cmult60} {iopath_Amult27_Cmult61} {iopath_Amult27_Cmult62} {iopath_Amult27_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult28_Cmult28} {iopath_Amult28_Cmult29} {iopath_Amult28_Cmult30} {iopath_Amult28_Cmult31} {iopath_Amult28_Cmult32} {iopath_Amult28_Cmult33} {iopath_Amult28_Cmult34} {iopath_Amult28_Cmult35} {iopath_Amult28_Cmult36} {iopath_Amult28_Cmult37} {iopath_Amult28_Cmult38} {iopath_Amult28_Cmult39} {iopath_Amult28_Cmult40} {iopath_Amult28_Cmult41} {iopath_Amult28_Cmult42} {iopath_Amult28_Cmult43} {iopath_Amult28_Cmult44} {iopath_Amult28_Cmult45} {iopath_Amult28_Cmult46} {iopath_Amult28_Cmult47} {iopath_Amult28_Cmult48} {iopath_Amult28_Cmult49} {iopath_Amult28_Cmult50} {iopath_Amult28_Cmult51} {iopath_Amult28_Cmult52} {iopath_Amult28_Cmult53} {iopath_Amult28_Cmult54} {iopath_Amult28_Cmult55} {iopath_Amult28_Cmult56} {iopath_Amult28_Cmult57} {iopath_Amult28_Cmult58} {iopath_Amult28_Cmult59} {iopath_Amult28_Cmult60} {iopath_Amult28_Cmult61} {iopath_Amult28_Cmult62} {iopath_Amult28_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult29_Cmult29} {iopath_Amult29_Cmult30} {iopath_Amult29_Cmult31} {iopath_Amult29_Cmult32} {iopath_Amult29_Cmult33} {iopath_Amult29_Cmult34} {iopath_Amult29_Cmult35} {iopath_Amult29_Cmult36} {iopath_Amult29_Cmult37} {iopath_Amult29_Cmult38} {iopath_Amult29_Cmult39} {iopath_Amult29_Cmult40} {iopath_Amult29_Cmult41} {iopath_Amult29_Cmult42} {iopath_Amult29_Cmult43} {iopath_Amult29_Cmult44} {iopath_Amult29_Cmult45} {iopath_Amult29_Cmult46} {iopath_Amult29_Cmult47} {iopath_Amult29_Cmult48} {iopath_Amult29_Cmult49} {iopath_Amult29_Cmult50} {iopath_Amult29_Cmult51} {iopath_Amult29_Cmult52} {iopath_Amult29_Cmult53} {iopath_Amult29_Cmult54} {iopath_Amult29_Cmult55} {iopath_Amult29_Cmult56} {iopath_Amult29_Cmult57} {iopath_Amult29_Cmult58} {iopath_Amult29_Cmult59} {iopath_Amult29_Cmult60} {iopath_Amult29_Cmult61} {iopath_Amult29_Cmult62} {iopath_Amult29_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult30_Cmult30} {iopath_Amult30_Cmult31} {iopath_Amult30_Cmult32} {iopath_Amult30_Cmult33} {iopath_Amult30_Cmult34} {iopath_Amult30_Cmult35} {iopath_Amult30_Cmult36} {iopath_Amult30_Cmult37} {iopath_Amult30_Cmult38} {iopath_Amult30_Cmult39} {iopath_Amult30_Cmult40} {iopath_Amult30_Cmult41} {iopath_Amult30_Cmult42} {iopath_Amult30_Cmult43} {iopath_Amult30_Cmult44} {iopath_Amult30_Cmult45} {iopath_Amult30_Cmult46} {iopath_Amult30_Cmult47} {iopath_Amult30_Cmult48} {iopath_Amult30_Cmult49} {iopath_Amult30_Cmult50} {iopath_Amult30_Cmult51} {iopath_Amult30_Cmult52} {iopath_Amult30_Cmult53} {iopath_Amult30_Cmult54} {iopath_Amult30_Cmult55} {iopath_Amult30_Cmult56} {iopath_Amult30_Cmult57} {iopath_Amult30_Cmult58} {iopath_Amult30_Cmult59} {iopath_Amult30_Cmult60} {iopath_Amult30_Cmult61} {iopath_Amult30_Cmult62} {iopath_Amult30_Cmult63} 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 0 {iopath_Amult31_Cmult31} {iopath_Amult31_Cmult32} {iopath_Amult31_Cmult33} {iopath_Amult31_Cmult34} {iopath_Amult31_Cmult35} {iopath_Amult31_Cmult36} {iopath_Amult31_Cmult37} {iopath_Amult31_Cmult38} {iopath_Amult31_Cmult39} {iopath_Amult31_Cmult40} {iopath_Amult31_Cmult41} {iopath_Amult31_Cmult42} {iopath_Amult31_Cmult43} {iopath_Amult31_Cmult44} {iopath_Amult31_Cmult45} {iopath_Amult31_Cmult46} {iopath_Amult31_Cmult47} {iopath_Amult31_Cmult48} {iopath_Amult31_Cmult49} {iopath_Amult31_Cmult50} {iopath_Amult31_Cmult51} {iopath_Amult31_Cmult52} {iopath_Amult31_Cmult53} {iopath_Amult31_Cmult54} {iopath_Amult31_Cmult55} {iopath_Amult31_Cmult56} {iopath_Amult31_Cmult57} {iopath_Amult31_Cmult58} {iopath_Amult31_Cmult59} {iopath_Amult31_Cmult60} {iopath_Amult31_Cmult61} {iopath_Amult31_Cmult62} {iopath_Amult31_Cmult63} "*)
	(* DELAY_MATRIX_Valid_mult="1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 "*)
	(* DELAY_MATRIX_sel_mul_32x32="1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 1e-10 "*)
	reg [63:0] Cmult_r;
	
    specify
		(Amult *> Cmult) = "";
		(Bmult *> Cmult) = "";
    endspecify
	
	assign Cmult = Cmult_r;
	
	always @(*) begin
		if (sel_mul_32x32 == 1'b1) begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult_r <= Amult * Bmult;
			end
		end else begin
			if (Valid_mult[0] == 1'b1) begin
				Cmult_r[31:0] <= Amult[15:0] * Bmult[15:0];
			end
			if (Valid_mult[1] == 1'b1) begin
				Cmult_r[63:32] <= Amult[31:16] * Bmult[31:16];
			end
		end
	end


endmodule
