`timescale 1ns / 10ps

module top (
    output wire [3:0] led
);

wire pwm0;
wire pwm1;
wire pwm2;

wire WB_CLK;
wire Clk_C16;
wire Clk_C16_Rst;
wire Clk_C21;
wire Clk_C21_Rst;
wire RST_FB21; 
wire CLK_FB21;

// Wishbone Bus Signals
//
wire    [16:0]  WBs_ADR        ; // Wishbone Address Bus
wire            WBs_CYC        ; // Wishbone Client Cycle  Strobe (i.e. Chip Select)
wire     [3:0]  WBs_BYTE_STB   ; // Wishbone Byte   Enables
wire            WBs_WE         ; // Wishbone Write  Enable Strobe
wire            WBs_RD         ; // Wishbone Read   Enable Strobe
wire            WBs_STB        ; // Wishbone Transfer      Strobe
wire    [31:0]  WBs_RD_DAT     ; // Wishbone Read   Data Bus
wire    [31:0]  WBs_WR_DAT     ; // Wishbone Write  Data Bus
wire            WBs_ACK        ; // Wishbone Client Acknowledge
wire     [1:0]  WBs_BTE        ; // Wishbone Client Burst Type Extension
wire     [2:0]  WBs_CTI        ; // Wishbone Client Cycle Type Identifier
wire            WB_RST         ; // Wishbone FPGA Reset
wire            WB_RST_FPGA    ; // Wishbone FPGA Reset
wire            WBs_ERR        ;

// Device ID
//
reg [31:0] Device_ID = 32'h0;

assign WBs_BTE = 2'h0;
assign WBs_CTI = 3'h0;

gclkbuff u_gclkbuff_reset ( .A(Clk_C16_Rst | WB_RST) , .Z(WB_RST_FPGA)   );
gclkbuff u_gclkbuff_clock ( .A(Clk_C16             ) , .Z(WB_CLK     )   ); // Clock 16

gclkbuff u_gclkbuff_reset1 ( .A(Clk_C21_Rst) , .Z(RST_FB21) );  
gclkbuff u_gclkbuff_clock1 ( .A(Clk_C21    ) , .Z(CLK_FB21) );  // Clock 21 

litex_core u_soc (
    .wb_adr ( WBs_ADR[16:2] ),
    .wb_dat_w ( WBs_WR_DAT ),
    .wb_dat_r ( WBs_RD_DAT ),
    .wb_sel ( WBs_BYTE_STB ),
    .wb_cyc ( WBs_CYC ),
    .wb_stb ( WBs_STB ),
    .wb_ack ( WBs_ACK ),
    .wb_we  ( WBs_WE  ),
    .wb_cti ( WBs_CTI ),
    .wb_bte ( WBs_BTE ),
    .sys_clk ( WB_CLK ),
    .wb_err ( WBs_ERR ),
    .pwm0( pwm0 ),
    .pwm0( pwm1 ),
    .pwm0( pwm2 ),
    .sys_rst ( WB_RST_FPGA ),
    );

// Empty Verilog model of QLAL4S3B
//
qlal4s3b_cell_macro              u_qlal4s3b_cell_macro
                               (
    // AHB-To-FPGA Bridge
    //
    .WBs_ADR                   ( WBs_ADR                     ), // output [16:0] | Address Bus                to   FPGA
    .WBs_CYC                   ( WBs_CYC                     ), // output        | Cycle Chip Select          to   FPGA
    .WBs_BYTE_STB              ( WBs_BYTE_STB                ), // output  [3:0] | Byte Select                to   FPGA
    .WBs_WE                    ( WBs_WE                      ), // output        | Write Enable               to   FPGA
    .WBs_RD                    ( WBs_RD                      ), // output        | Read  Enable               to   FPGA
    .WBs_STB                   ( WBs_STB                     ), // output        | Strobe Signal              to   FPGA
    .WBs_WR_DAT                ( WBs_WR_DAT                  ), // output [31:0] | Write Data Bus             to   FPGA
    .WB_CLK                    ( WB_CLK                      ), // input         | FPGA Clock               from FPGA
    .WB_RST                    ( WB_RST                      ), // output        | FPGA Reset               to   FPGA
    .WBs_RD_DAT                ( WBs_RD_DAT                  ), // input  [31:0] | Read Data Bus              from FPGA
    .WBs_ACK                   ( WBs_ACK                     ), // input         | Transfer Cycle Acknowledge from FPGA
    //
    // SDMA Signals
    //
    .SDMA_Req                  (  4'h0  					 ), // input   [3:0]
    .SDMA_Sreq                 (  4'h0                       ), // input   [3:0]
    .SDMA_Done                 (							 ), // output  [3:0]
    .SDMA_Active               (							 ), // output  [3:0]
    //
    // FB Interrupts
    //
    .FB_msg_out                (  4'h0                       ), // input   [3:0]
    .FB_Int_Clr                (  8'h0                       ), // input   [7:0]
    .FB_Start                  (                             ), // output
    .FB_Busy                   (  1'b0                       ), // input
    //
    // FB Clocks
    //
    .Clk_C16                   ( Clk_C16                     ), // output
    .Clk_C16_Rst               ( Clk_C16_Rst                 ), // output
    .Clk_C21                   ( Clk_C21                     ), // output
    .Clk_C21_Rst               ( Clk_C21_Rst                 ), // output
    //
    // Packet FIFO
    //
    .Sys_PKfb_Clk              (  1'b0                       ), // input
    .Sys_PKfb_Rst              (                             ), // output
    .FB_PKfbData               ( 32'h0                       ), // input  [31:0]
    .FB_PKfbPush               (  4'h0                       ), // input   [3:0]
    .FB_PKfbSOF                (  1'b0                       ), // input
    .FB_PKfbEOF                (  1'b0                       ), // input
    .FB_PKfbOverflow           (                             ), // output
	//
	// Sensor Interface
	//
    .Sensor_Int                (                             ), // output  [7:0]
    .TimeStamp                 (                             ), // output [23:0]
    //
    // SPI Master APB Bus
    //
    .Sys_Pclk                  (                             ), // output
    .Sys_Pclk_Rst              (                             ), // output      <-- Fixed to add "_Rst"
    .Sys_PSel                  (  1'b0                       ), // input
    .SPIm_Paddr                ( 16'h0                       ), // input  [15:0]
    .SPIm_PEnable              (  1'b0                       ), // input
    .SPIm_PWrite               (  1'b0                       ), // input
    .SPIm_PWdata               ( 32'h0                       ), // input  [31:0]
    .SPIm_Prdata               (                             ), // output [31:0]
    .SPIm_PReady               (                             ), // output
    .SPIm_PSlvErr              (                             ), // output
    //
    // Misc
    //
    .Device_ID                 ( Device_ID[19:4]             ), // input  [15:0]
    //
    // FBIO Signals
    //
    .FBIO_In                   (                             ), // output [13:0] <-- Do Not make any connections; Use Constraint manager in SpDE to sFBIO
    .FBIO_In_En                (                             ), // input  [13:0] <-- Do Not make any connections; Use Constraint manager in SpDE to sFBIO
    .FBIO_Out                  (                             ), // input  [13:0] <-- Do Not make any connections; Use Constraint manager in SpDE to sFBIO
    .FBIO_Out_En               (                             ), // input  [13:0] <-- Do Not make any connections; Use Constraint manager in SpDE to sFBIO
	//
	// ???
	//
    .SFBIO                     (                             ), // inout  [13:0]
    .Device_ID_6S              ( 1'b0                        ), // input
    .Device_ID_4S              ( 1'b0                        ), // input
    .SPIm_PWdata_26S           ( 1'b0                        ), // input
    .SPIm_PWdata_24S           ( 1'b0                        ), // input
    .SPIm_PWdata_14S           ( 1'b0                        ), // input
    .SPIm_PWdata_11S           ( 1'b0                        ), // input
    .SPIm_PWdata_0S            ( 1'b0                        ), // input
    .SPIm_Paddr_8S             ( 1'b0                        ), // input
    .SPIm_Paddr_6S             ( 1'b0                        ), // input
    .FB_PKfbPush_1S            ( 1'b0                        ), // input
    .FB_PKfbData_31S           ( 1'b0                        ), // input
    .FB_PKfbData_21S           ( 1'b0                        ), // input
    .FB_PKfbData_19S           ( 1'b0                        ), // input
    .FB_PKfbData_9S            ( 1'b0                        ), // input
    .FB_PKfbData_6S            ( 1'b0                        ), // input
    .Sys_PKfb_ClkS             ( 1'b0                        ), // input
    .FB_BusyS                  ( 1'b0                        ), // input
    .WB_CLKS                   ( 1'b0                        )  // input
                                                             );

// ============================================================================

// A counter for blinking led
reg [19:0] cnt;
initial cnt <= 0;

always @(posedge WB_CLK)
    if (WB_RST_FPGA)
        cnt <= 0;
    else
        cnt <= cnt + 1;

// LED connections
assign led[0] = pwm0;
assign led[2] = pwm1;
assign led[1] = pwm2;
assign led[3] = cnt[19];

endmodule
